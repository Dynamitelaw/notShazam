`define NFFT 256 // if change this, change FREQ_WIDTH
`define FREQS (`NFFT / 2)
`define FREQ_WIDTH 7 // if change NFFT, change this

`define FINAL_AMPL_WIDTH 24
`define INPUT_AMPL_WIDTH 24

`define PEAKS 6 // Changing this requires many changes in code
