// CSEE 4840 Design Project
// By: Jose Rubianes & Tomin Perea-Chamblee & Eitan Kaplan


`include "./AudioCodecDrivers/audio_driver.sv"
//`include "SfftPipeline.sv"
`include "SfftPipeline_SingleStage.sv"
//`include "peaks.sv"
//`include "peaksSequential.sv"


module FFT_Accelerator( 
		  input logic clk,
		  input logic reset,

		  input logic [3:0] 	KEY, // Pushbuttons; KEY[0] is rightmost

		  // 7-segment LED displays; HEX0 is rightmost
		  output logic [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5,
		  
		  //Audio pin assignments
		  output logic FPGA_I2C_SCLK,
		  inout FPGA_I2C_SDAT,
		  output logic AUD_XCK,
		  input logic AUD_DACLRCK,
		  input logic AUD_ADCLRCK,
		  input logic AUD_BCLK,
		  input logic AUD_ADCDAT,
		  output logic AUD_DACDAT,
		  
		  //Driver IO ports
		  input logic [7:0] writedata,
		  input logic write,
		  input chipselect,
		  input logic [15:0] address,
		  output logic [7:0] readdata
		  );

	
	/*
	//Debounce button inputs 
	wire KEY3db, KEY2db, KEY1db, KEY0db;  //debounced buttons
	debouncer db(.clk(clk), .buttonsIn(KEY), .buttonsOut({KEY3db, KEY2db, KEY1db, KEY0db}));
	*/
	
	//Instantiate audio controller
	reg [23:0] dac_left_in;
	reg [23:0] dac_right_in;
	
	wire [23:0] adc_left_out;
	wire [23:0] adc_right_out;
	
	wire advance;
	
	reg [23:0] adc_out_buffer = 0;
	
	reg [24:0] counter = 0;  //downsample adance signal
	
	audio_driver aDriver(
	 	.CLOCK_50(clk), 
	 	.reset(reset), 
	 	.dac_left(dac_left_in), 
	 	.dac_right(dac_right_in), 
	 	.adc_left(adc_left_out), 
	 	.adc_right(adc_right_out), 
	 	.advance(advance), 
	 	.FPGA_I2C_SCLK(FPGA_I2C_SCLK), 
	 	.FPGA_I2C_SDAT(FPGA_I2C_SDAT), 
	 	.AUD_XCK(AUD_XCK), 
	 	.AUD_DACLRCK(AUD_DACLRCK), 
	 	.AUD_ADCLRCK(AUD_ADCLRCK), 
	 	.AUD_BCLK(AUD_BCLK), 
	 	.AUD_ADCDAT(AUD_ADCDAT), 
	 	.AUD_DACDAT(AUD_DACDAT)
	 	);
	 
	//Convert stereo input to mono	
	//500 Hz test wave
	reg [23:0] testWave [43999:0] = '{24'd8388608, 
24'd8706954, 24'd8962301, 24'd9104115, 24'd9104331, 24'd8962907, 24'd8707830, 24'd8389579, 24'd8071136, 24'd7815521, 24'd7673317, 24'd7672669, 24'd7813703, 24'd8068510, 24'd8386664, 24'd8705202, 24'd8961087, 24'd9103679, 24'd9104760, 24'd8964115, 24'd8709579, 24'd8391523, 24'd8072890, 24'd7816737, 24'd7673756, 24'd7672243, 24'd7812497, 24'd8066762, 24'd8384720, 24'd8703447, 24'd8959868, 
24'd9103238, 24'd9105183, 24'd8965320, 24'd8711326, 24'd8393466, 24'd8074646, 24'd7817957, 24'd7674200, 24'd7671822, 24'd7811295, 24'd8065017, 24'd8382777, 24'd8701691, 24'd8958646, 24'd9102792, 24'd9105602, 24'd8966520, 24'd8713070, 24'd8395410, 24'd8076404, 24'd7819182, 24'd7674648, 24'd7671406, 24'd7810097, 24'd8063273, 24'd8380833, 24'd8699932, 24'd8957420, 24'd9102341, 24'd9106015, 
24'd8967716, 24'd8714812, 24'd8397353, 24'd8078164, 24'd7820410, 24'd7675102, 24'd7670995, 24'd7808902, 24'd8061532, 24'd8378890, 24'd8698171, 24'd8956189, 24'd9101884, 24'd9106424, 24'd8968908, 24'd8716552, 24'd8399297, 24'd8079926, 24'd7821643, 24'd7675560, 24'd7670589, 24'd7807712, 24'd8059794, 24'd8376947, 24'd8696407, 24'd8954955, 24'd9101423, 24'd9106827, 24'd8970096, 24'd8718290, 
24'd8401240, 24'd8081690, 24'd7822879, 24'd7676024, 24'd7670188, 24'd7806526, 24'd8058057, 24'd8375003, 24'd8694642, 24'd8953716, 24'd9100957, 24'd9107225, 24'd8971280, 24'd8720025, 24'd8403183, 24'd8083457, 24'd7824119, 24'd7676493, 24'd7669792, 24'd7805344, 24'd8056323, 24'd8373060, 24'd8692874, 24'd8952474, 24'd9100486, 24'd9107619, 24'd8972460, 24'd8721758, 24'd8405127, 24'd8085226, 
24'd7825363, 24'd7676966, 24'd7669402, 24'd7804166, 24'd8054591, 24'd8371117, 24'd8691104, 24'd8951228, 24'd9100010, 24'd9108007, 24'd8973636, 24'd8723489, 24'd8407070, 24'd8086996, 24'd7826612, 24'd7677445, 24'd7669016, 24'd7802993, 24'd8052862, 24'd8369174, 24'd8689332, 24'd8949978, 24'd9099529, 24'd9108390, 24'd8974808, 24'd8725217, 24'd8409012, 24'd8088769, 24'd7827864, 24'd7677928, 
24'd7668635, 24'd7801823, 24'd8051134, 24'd8367231, 24'd8687558, 24'd8948724, 24'd9099043, 24'd9108768, 24'd8975975, 24'd8726943, 24'd8410955, 24'd8090545, 24'd7829120, 24'd7678417, 24'd7668259, 24'd7800657, 24'd8049410, 24'd8365288, 24'd8685782, 24'd8947466, 24'd9098552, 24'd9109142, 24'd8977139, 24'd8728667, 24'd8412898, 24'd8092322, 24'd7830380, 24'd7678911, 24'd7667889, 24'd7799496, 
24'd8047687, 24'd8363346, 24'd8684004, 24'd8946204, 24'd9098056, 24'd9109510, 24'd8978298, 24'd8730388, 24'd8414840, 24'd8094101, 24'd7831644, 24'd7679409, 24'd7667523, 24'd7798339, 24'd8045967, 24'd8361404, 24'd8682224, 24'd8944938, 24'd9097555, 24'd9109873, 24'd8979453, 24'd8732107, 24'd8416782, 24'd8095882, 24'd7832912, 24'd7679913, 24'd7667163, 24'd7797185, 24'd8044250, 24'd8359461, 
24'd8680441, 24'd8943668, 24'd9097049, 24'd9110231, 24'd8980605, 24'd8733823, 24'd8418724, 24'd8097666, 24'd7834184, 24'd7680421, 24'd7666807, 24'd7796036, 24'd8042534, 24'd8357520, 24'd8678657, 24'd8942394, 24'd9096538, 24'd9110584, 24'd8981752, 24'd8735537, 24'd8420666, 24'd8099451, 24'd7835459, 24'd7680934, 24'd7666457, 24'd7794892, 24'd8040822, 24'd8355578, 24'd8676871, 24'd8941117, 
24'd9096022, 24'd9110931, 24'd8982894, 24'd8737249, 24'd8422608, 24'd8101238, 24'd7836739, 24'd7681453, 24'd7666111, 24'd7793751, 24'd8039111, 24'd8353636, 24'd8675082, 24'd8939835, 24'd9095501, 24'd9111274, 24'd8984033, 24'd8738958, 24'd8424549, 24'd8103028, 24'd7838022, 24'd7681976, 24'd7665771, 24'd7792614, 24'd8037403, 24'd8351695, 24'd8673292, 24'd8938550, 24'd9094975, 24'd9111612, 
24'd8985167, 24'd8740665, 24'd8426490, 24'd8104819, 24'd7839309, 24'd7682504, 24'd7665436, 24'd7791482, 24'd8035698, 24'd8349754, 24'd8671499, 24'd8937261, 24'd9094445, 24'd9111945, 24'd8986298, 24'd8742369, 24'd8428431, 24'd8106613, 24'd7840600, 24'd7683038, 24'd7665106, 24'd7790354, 24'd8033995, 24'd8347813, 24'd8669705, 24'd8935968, 24'd9093909, 24'd9112272, 24'd8987424, 24'd8744071, 
24'd8430372, 24'd8108408, 24'd7841895, 24'd7683576, 24'd7664781, 24'd7789230, 24'd8032295, 24'd8345873, 24'd8667908, 24'd8934671, 24'd9093368, 24'd9112595, 24'd8988546, 24'd8745770, 24'd8432312, 24'd8110205, 24'd7843194, 24'd7684119, 24'd7664461, 24'd7788110, 24'd8030597, 24'd8343933, 24'd8666110, 24'd8933370, 24'd9092823, 24'd9112912, 24'd8989663, 24'd8747466, 24'd8434252, 24'd8112005, 
24'd7844497, 24'd7684667, 24'd7664146, 24'd7786994, 24'd8028901, 24'd8341993, 24'd8664310, 24'd8932066, 24'd9092272, 24'd9113225, 24'd8990777, 24'd8749161, 24'd8436192, 24'd8113806, 24'd7845803, 24'd7685220, 24'd7663836, 24'd7785883, 24'd8027208, 24'd8340054, 24'd8662508, 24'd8930757, 24'd9091717, 24'd9113532, 24'd8991886, 24'd8750852, 24'd8438131, 24'd8115609, 24'd7847113, 24'd7685778, 
24'd7663531, 24'd7784776, 24'd8025518, 24'd8338114, 24'd8660703, 24'd8929445, 24'd9091156, 24'd9113834, 24'd8992991, 24'd8752541, 24'd8440070, 24'd8117414, 24'd7848427, 24'd7686341, 24'd7663232, 24'd7783673, 24'd8023830, 24'd8336176, 24'd8658897, 24'd8928129, 24'd9090591, 24'd9114131, 24'd8994092, 24'd8754228, 24'd8442009, 24'd8119221, 24'd7849745, 24'd7686909, 24'd7662937, 24'd7782574, 
24'd8022145, 24'd8334237, 24'd8657089, 24'd8926810, 24'd9090021, 24'd9114423, 24'd8995188, 24'd8755912, 24'd8443947, 24'd8121030, 24'd7851067, 24'd7687481, 24'd7662648, 24'd7781480, 24'd8020462, 24'd8332299, 24'd8655280, 24'd8925486, 24'd9089445, 24'd9114710, 24'd8996281, 24'd8757593, 24'd8445885, 24'd8122841, 24'd7852392, 24'd7688059, 24'd7662363, 24'd7780390, 24'd8018782, 24'd8330361, 
24'd8653468, 24'd8924159, 24'd9088865, 24'd9114992, 24'd8997369, 24'd8759272, 24'd8447822, 24'd8124654, 24'd7853721, 24'd7688641, 24'd7662084, 24'd7779304, 24'd8017104, 24'd8328424, 24'd8651654, 24'd8922828, 24'd9088280, 24'd9115269, 24'd8998452, 24'd8760949, 24'd8449759, 24'd8126468, 24'd7855054, 24'd7689229, 24'd7661810, 24'd7778222, 24'd8015429, 24'd8326487, 24'd8649839, 24'd8921493, 
24'd9087690, 24'd9115540, 24'd8999532, 24'd8762622, 24'd8451696, 24'd8128284, 24'd7856390, 24'd7689821, 24'd7661541, 24'd7777145, 24'd8013757, 24'd8324551, 24'd8648022, 24'd8920155, 24'd9087096, 24'd9115807, 24'd9000607, 24'd8764293, 24'd8453632, 24'd8130103, 24'd7857731, 24'd7690419, 24'd7661277, 24'd7776072, 24'd8012087, 24'd8322615, 24'd8646203, 24'd8918813, 24'd9086496, 24'd9116068, 
24'd9001678, 24'd8765962, 24'd8455568, 24'd8131923, 24'd7859075, 24'd7691021, 24'd7661018, 24'd7775003, 24'd8010420, 24'd8320680, 24'd8644382, 24'd8917467, 24'd9085891, 24'd9116325, 24'd9002744, 24'd8767627, 24'd8457503, 24'd8133744, 24'd7860423, 24'd7691628, 24'd7660764, 24'd7773939, 24'd8008756, 24'd8318745, 24'd8642559, 24'd8916117, 24'd9085282, 24'd9116576, 24'd9003807, 24'd8769290, 
24'd8459438, 24'd8135568, 24'd7861774, 24'd7692240, 24'd7660515, 24'd7772879, 24'd8007094, 24'd8316810, 24'd8640735, 24'd8914764, 24'd9084668, 24'd9116822, 24'd9004865, 24'd8770951, 24'd8461372, 24'd8137393, 24'd7863129, 24'd7692856, 24'd7660272, 24'd7771823, 24'd8005435, 24'd8314876, 24'd8638909, 24'd8913407, 24'd9084048, 24'd9117063, 24'd9005918, 24'd8772609, 24'd8463306, 24'd8139220, 
24'd7864488, 24'd7693478, 24'd7660033, 24'd7770772, 24'd8003779, 24'd8312943, 24'd8637081, 24'd8912046, 24'd9083424, 24'd9117299, 24'd9006968, 24'd8774264, 24'd8465239, 24'd8141049, 24'd7865851, 24'd7694105, 24'd7659800, 24'd7769724, 24'd8002125, 24'd8311010, 24'd8635251, 24'd8910682, 24'd9082795, 24'd9117530, 24'd9008013, 24'd8775916, 24'd8467172, 24'd8142880, 24'd7867217, 24'd7694736, 
24'd7659571, 24'd7768682, 24'd8000474, 24'd8309077, 24'd8633419, 24'd8909314, 24'd9082161, 24'd9117756, 24'd9009053, 24'd8777566, 24'd8469104, 24'd8144712, 24'd7868587, 24'd7695372, 24'd7659348, 24'd7767643, 24'd7998826, 24'd8307145, 24'd8631586, 24'd8907942, 24'd9081523, 24'd9117976, 24'd9010090, 24'd8779212, 24'd8471035, 24'd8146546, 24'd7869960, 24'd7696014, 24'd7659130, 24'd7766609, 
24'd7997180, 24'd8305214, 24'd8629751, 24'd8906567, 24'd9080879, 24'd9118192, 24'd9011121, 24'd8780857, 24'd8472966, 24'd8148382, 24'd7871337, 24'd7696660, 24'd7658917, 24'd7765579, 24'd7995537, 24'd8303283, 24'd8627915, 24'd8905188, 24'd9080231, 24'd9118402, 24'd9012149, 24'd8782498, 24'd8474897, 24'd8150219, 24'd7872718, 24'd7697310, 24'd7658709, 24'd7764554, 24'd7993897, 24'd8301353, 
24'd8626077, 24'd8903805, 24'd9079577, 24'd9118608, 24'd9013172, 24'd8784137, 24'd8476827, 24'd8152058, 24'd7874102, 24'd7697966, 24'd7658507, 24'd7763533, 24'd7992260, 24'd8299424, 24'd8624237, 24'd8902419, 24'd9078919, 24'd9118808, 24'd9014191, 24'd8785772, 24'd8478756, 24'd8153899, 24'd7875490, 24'd7698627, 24'd7658309, 24'd7762516, 24'd7990626, 24'd8297495, 24'd8622395, 24'd8901029, 
24'd9078256, 24'd9119003, 24'd9015205, 24'd8787406, 24'd8480684, 24'd8155741, 24'd7876882, 24'd7699292, 24'd7658117, 24'd7761504, 24'd7988994, 24'd8295567, 24'd8620552, 24'd8899636, 24'd9077588, 24'd9119193, 24'd9016216, 24'd8789036, 24'd8482612, 24'd8157585, 24'd7878277, 24'd7699962, 24'd7657929, 24'd7760496, 24'd7987365, 24'd8293639, 24'd8618707, 24'd8898239, 24'd9076916, 24'd9119377, 
24'd9017221, 24'd8790663, 24'd8484539, 24'd8159431, 24'd7879676, 24'd7700637, 24'd7657747, 24'd7759493, 24'd7985739, 24'd8291712, 24'd8616861, 24'd8896839, 24'd9076238, 24'd9119557, 24'd9018222, 24'd8792288, 24'd8486466, 24'd8161278, 24'd7881078, 24'd7701317, 24'd7657570, 24'd7758494, 24'd7984116, 24'd8289786, 24'd8615013, 24'd8895435, 24'd9075556, 24'd9119732, 24'd9019219, 24'd8793910, 
24'd8488392, 24'd8163127, 24'd7882484, 24'd7702002, 24'd7657398, 24'd7757499, 24'd7982495, 24'd8287861, 24'd8613163, 24'd8894027, 24'd9074869, 24'd9119901, 24'd9020212, 24'd8795529, 24'd8490317, 24'd8164977, 24'd7883893, 24'd7702691, 24'd7657231, 24'd7756509, 24'd7980878, 24'd8285936, 24'd8611312, 24'd8892616, 24'd9074177, 24'd9120065, 24'd9021200, 24'd8797145, 24'd8492241, 24'd8166829, 
24'd7885306, 24'd7703386, 24'd7657069, 24'd7755523, 24'd7979263, 24'd8284012, 24'd8609459, 24'd8891201, 24'd9073480, 24'd9120225, 24'd9022183, 24'd8798758, 24'd8494165, 24'd8168683, 24'd7886723, 24'd7704085, 24'd7656913, 24'd7754542, 24'd7977651, 24'd8282088, 24'd8607605, 24'd8889783, 24'd9072779, 24'd9120379, 24'd9023162, 24'd8800369, 24'd8496088, 24'd8170538, 24'd7888143, 24'd7704789, 
24'd7656761, 24'd7753565, 24'd7976042, 24'd8280166, 24'd8605749, 24'd8888361, 24'd9072072, 24'd9120527, 24'd9024137, 24'd8801976, 24'd8498010, 24'd8172394, 24'd7889566, 24'd7705497, 24'd7656615, 24'd7752593, 24'd7974436, 24'd8278244, 24'd8603892, 24'd8886936, 24'd9071361, 24'd9120671, 24'd9025107, 24'd8803581, 24'd8499932, 24'd8174252, 24'd7890993, 24'd7706211, 24'd7656474, 24'd7751625, 
24'd7972833, 24'd8276323, 24'd8602033, 24'd8885507, 24'd9070645, 24'd9120810, 24'd9026073, 24'd8805182, 24'd8501853, 24'd8176112, 24'd7892424, 24'd7706929, 24'd7656338, 24'd7750661, 24'd7971233, 24'd8274402, 24'd8600173, 24'd8884075, 24'd9069925, 24'd9120943, 24'd9027034, 24'd8806781, 24'd8503773, 24'd8177973, 24'd7893858, 24'd7707652, 24'd7656207, 24'd7749702, 24'd7969636, 24'd8272483, 
24'd8598311, 24'd8882639, 24'd9069199, 24'd9121072, 24'd9027991, 24'd8808377, 24'd8505692, 24'd8179836, 24'd7895295, 24'd7708380, 24'd7656081, 24'd7748748, 24'd7968041, 24'd8270564, 24'd8596448, 24'd8881200, 24'd9068469, 24'd9121195, 24'd9028943, 24'd8809970, 24'd8507610, 24'd8181700, 24'd7896736, 24'd7709113, 24'd7655960, 24'd7747798, 24'd7966450, 24'd8268646, 24'd8594583, 24'd8879757, 
24'd9067734, 24'd9121313, 24'd9029891, 24'd8811560, 24'd8509527, 24'd8183565, 24'd7898180, 24'd7709850, 24'd7655845, 24'd7746852, 24'd7964861, 24'd8266729, 24'd8592717, 24'd8878311, 24'd9066994, 24'd9121426, 24'd9030834, 24'd8813147, 24'd8511444, 24'd8185432, 24'd7899628, 24'd7710592, 24'd7655734, 24'd7745911, 24'd7963276, 24'd8264813, 24'd8590849, 24'd8876862, 24'd9066250, 24'd9121534, 
24'd9031773, 24'd8814731, 24'd8513360, 24'd8187300, 24'd7901079, 24'd7711339, 24'd7655629, 24'd7744974, 24'd7961693, 24'd8262898, 24'd8588980, 24'd8875409, 24'd9065501, 24'd9121636, 24'd9032707, 24'd8816312, 24'd8515275, 24'd8189170, 24'd7902534, 24'd7712091, 24'd7655529, 24'd7744042, 24'd7960114, 24'd8260983, 24'd8587110, 24'd8873952, 24'd9064747, 24'd9121734, 24'd9033637, 24'd8817890, 
24'd8517189, 24'd8191041, 24'd7903992, 24'd7712847, 24'd7655434, 24'd7743115, 24'd7958537, 24'd8259070, 24'd8585238, 24'd8872493, 24'd9063988, 24'd9121826, 24'd9034562, 24'd8819465, 24'd8519102, 24'd8192914, 24'd7905453, 24'd7713608, 24'd7655344, 24'd7742192, 24'd7956964, 24'd8257157, 24'd8583364, 24'd8871030, 24'd9063224, 24'd9121914, 24'd9035483, 24'd8821037, 24'd8521014, 24'd8194788, 
24'd7906918, 24'd7714374, 24'd7655260, 24'd7741273, 24'd7955393, 24'd8255246, 24'd8581490, 24'd8869563, 24'd9062456, 24'd9121996, 24'd9036399, 24'd8822606, 24'd8522925, 24'd8196663, 24'd7908386, 24'd7715145, 24'd7655180, 24'd7740359, 24'd7953826, 24'd8253335, 24'd8579614, 24'd8868093, 24'd9061683, 24'd9122073, 24'd9037311, 24'd8824172, 24'd8524835, 24'd8198540, 24'd7909858, 24'd7715920, 
24'd7655106, 24'd7739450, 24'd7952261, 24'd8251425, 24'd8577737, 24'd8866620, 24'd9060906, 24'd9122145, 24'd9038218, 24'd8825735, 24'd8526745, 24'd8200418, 24'd7911333, 24'd7716700, 24'd7655036, 24'd7738545, 24'd7950700, 24'd8249516, 24'd8575858, 24'd8865143, 24'd9060123, 24'd9122211, 24'd9039120, 24'd8827294, 24'd8528653, 24'd8202297, 24'd7912811, 24'd7717485, 24'd7654972, 24'd7737645, 
24'd7949142, 24'd8247608, 24'd8573978, 24'd8863663, 24'd9059336, 24'd9122273, 24'd9040018, 24'd8828851, 24'd8530560, 24'd8204177, 24'd7914293, 24'd7718274, 24'd7654913, 24'd7736749, 24'd7947587, 24'd8245701, 24'd8572097, 24'd8862180, 24'd9058544, 24'd9122329, 24'd9040912, 24'd8830405, 24'd8532467, 24'd8206059, 24'd7915778, 24'd7719068, 24'd7654860, 24'd7735858, 24'd7946035, 24'd8243795, 
24'd8570214, 24'd8860694, 24'd9057748, 24'd9122380, 24'd9041801, 24'd8831955, 24'd8534372, 24'd8207942, 24'd7917266, 24'd7719867, 24'd7654811, 24'd7734972, 24'd7944486, 24'd8241891, 24'd8568331, 24'd8859204, 24'd9056947, 24'd9122427, 24'd9042685, 24'd8833503, 24'd8536276, 24'd8209827, 24'd7918758, 24'd7720671, 24'd7654767, 24'd7734090, 24'd7942940, 24'd8239987, 24'd8566446, 24'd8857710, 
24'd9056141, 24'd9122468, 24'd9043565, 24'd8835047, 24'd8538180, 24'd8211712, 24'd7920252, 24'd7721479, 24'd7654729, 24'd7733212, 24'd7941397, 24'd8238084, 24'd8564559, 24'd8856214, 24'd9055330, 24'd9122503, 24'd9044440, 24'd8836588, 24'd8540082, 24'd8213599, 24'd7921751, 24'd7722292, 24'd7654696, 24'd7732339, 24'd7939857, 24'd8236182, 24'd8562672, 24'd8854714, 24'd9054515, 24'd9122534, 
24'd9045310, 24'd8838126, 24'd8541983, 24'd8215488, 24'd7923252, 24'd7723109, 24'd7654668, 24'd7731471, 24'd7938321, 24'd8234282, 24'd8560783, 24'd8853211, 24'd9053695, 24'd9122560, 24'd9046176, 24'd8839661, 24'd8543883, 24'd8217377, 24'd7924757, 24'd7723932, 24'd7654645, 24'd7730608, 24'd7936788, 24'd8232382, 24'd8558893, 24'd8851705, 24'd9052871, 24'd9122580, 24'd9047037, 24'd8841193, 
24'd8545782, 24'd8219267, 24'd7926265, 24'd7724758, 24'd7654627, 24'd7729749, 24'd7935258, 24'd8230483, 24'd8557002, 24'd8850195, 24'd9052041, 24'd9122595, 24'd9047894, 24'd8842721, 24'd8547680, 24'd8221159, 24'd7927776, 24'd7725590, 24'd7654614, 24'd7728894, 24'd7933731, 24'd8228586, 24'd8555110, 24'd8848683, 24'd9051208, 24'd9122605, 24'd9048746, 24'd8844247, 24'd8549577, 24'd8223052, 
24'd7929290, 24'd7726426, 24'd7654607, 24'd7728045, 24'd7932207, 24'd8226690, 24'd8553216, 24'd8847167, 24'd9050369, 24'd9122610, 24'd9049593, 24'd8845769, 24'd8551473, 24'd8224946, 24'd7930808, 24'd7727267, 24'd7654604, 24'd7727200, 24'd7930686, 24'd8224795, 24'd8551321, 24'd8845647, 24'd9049526, 24'd9122610, 24'd9050436, 24'd8847288, 24'd8553367, 24'd8226841, 24'd7932328, 24'd7728112, 
24'd7654607, 24'd7726359, 24'd7929169, 24'd8222901, 24'd8549426, 24'd8844125, 24'd9048678, 24'd9122605, 24'd9051274, 24'd8848804, 24'd8555261, 24'd8228738, 24'd7933853, 24'd7728962, 24'd7654615, 24'd7725523, 24'd7927655, 24'd8221008, 24'd8547529, 24'd8842599, 24'd9047826, 24'd9122594, 24'd9052108, 24'd8850316, 24'd8557153, 24'd8230635, 24'd7935380, 24'd7729817, 24'd7654628, 24'd7724692, 
24'd7926144, 24'd8219116, 24'd8545631, 24'd8841070, 24'd9046969, 24'd9122578, 24'd9052937, 24'd8851825, 24'd8559044, 24'd8232534, 24'd7936910, 24'd7730677, 24'd7654646, 24'd7723866, 24'd7924636, 24'd8217226, 24'd8543732, 24'd8839538, 24'd9046107, 24'd9122558, 24'd9053761, 24'd8853331, 24'd8560934, 24'd8234433, 24'd7938444, 24'd7731540, 24'd7654670, 24'd7723044, 24'd7923132, 24'd8215337, 
24'd8541831, 24'd8838003, 24'd9045241, 24'd9122532, 24'd9054580, 24'd8854834, 24'd8562823, 24'd8236334, 24'd7939980, 24'd7732409, 24'd7654698, 24'd7722227, 24'd7921631, 24'd8213448, 24'd8539930, 24'd8836465, 24'd9044370, 24'd9122501, 24'd9055395, 24'd8856334, 24'd8564710, 24'd8238236, 24'd7941520, 24'd7733282, 24'd7654732, 24'd7721414, 24'd7920133, 24'd8211562, 24'd8538028, 24'd8834924, 
24'd9043495, 24'd9122464, 24'd9056205, 24'd8857830, 24'd8566596, 24'd8240139, 24'd7943063, 24'd7734160, 24'd7654771, 24'd7720606, 24'd7918638, 24'd8209676, 24'd8536124, 24'd8833379, 24'd9042614, 24'd9122423, 24'd9057011, 24'd8859323, 24'd8568481, 24'd8242043, 24'd7944609, 24'd7735042, 24'd7654815, 24'd7719803, 24'd7917147, 24'd8207792, 24'd8534220, 24'd8831831, 24'd9041730, 24'd9122377, 
24'd9057812, 24'd8860813, 24'd8570365, 24'd8243948, 24'd7946159, 24'd7735929, 24'd7654864, 24'd7719005, 24'd7915659, 24'd8205909, 24'd8532314, 24'd8830281, 24'd9040841, 24'd9122325, 24'd9058608, 24'd8862299, 24'd8572247, 24'd8245854, 24'd7947711, 24'd7736821, 24'd7654918, 24'd7718211, 24'd7914174, 24'd8204027, 24'd8530408, 24'd8828727, 24'd9039947, 24'd9122268, 24'd9059399, 24'd8863782, 
24'd8574128, 24'd8247761, 24'd7949266, 24'd7737717, 24'd7654977, 24'd7717422, 24'd7912693, 24'd8202147, 24'd8528500, 24'd8827170, 24'd9039048, 24'd9122206, 24'd9060186, 24'd8865262, 24'd8576008, 24'd8249669, 24'd7950825, 24'd7738617, 24'd7655042, 24'd7716638, 24'd7911215, 24'd8200267, 24'd8526592, 24'd8825610, 24'd9038146, 24'd9122139, 24'd9060968, 24'd8866738, 24'd8577887, 24'd8251578, 
24'd7952386, 24'd7739523, 24'd7655111, 24'd7715858, 24'd7909740, 24'd8198390, 24'd8524683, 24'd8824047, 24'd9037238, 24'd9122067, 24'd9061745, 24'd8868211, 24'd8579764, 24'd8253487, 24'd7953951, 24'd7740432, 24'd7655186, 24'd7715083, 24'd7908269, 24'd8196513, 24'd8522772, 24'd8822480, 24'd9036326, 24'd9121989, 24'd9062518, 24'd8869680, 24'd8581640, 24'd8255398, 24'd7955519, 24'd7741347, 
24'd7655266, 24'd7714313, 24'd7906801, 24'd8194638, 24'd8520861, 24'd8820911, 24'd9035410, 24'd9121907, 24'd9063286, 24'd8871147, 24'd8583514, 24'd8257310, 24'd7957089, 24'd7742265, 24'd7655351, 24'd7713547, 24'd7905336, 24'd8192764, 24'd8518949, 24'd8819339, 24'd9034488, 24'd9121819, 24'd9064049, 24'd8872610, 24'd8585387, 24'd8259223, 24'd7958663, 24'd7743189, 24'd7655442, 24'd7712787, 
24'd7903875, 24'd8190892, 24'd8517036, 24'd8817764, 24'd9033563, 24'd9121726, 24'd9064807, 24'd8874069, 24'd8587259, 24'd8261136, 24'd7960240, 24'd7744117, 24'd7655537, 24'd7712031, 24'd7902417, 24'd8189021, 24'd8515122, 24'd8816186, 24'd9032633, 24'd9121628, 24'd9065561, 24'd8875525, 24'd8589129, 24'd8263051, 24'd7961820, 24'd7745049, 24'd7655637, 24'd7711279, 24'd7900963, 24'd8187151, 
24'd8513207, 24'd8814604, 24'd9031698, 24'd9121525, 24'd9066310, 24'd8876978, 24'd8590998, 24'd8264966, 24'd7963402, 24'd7745986, 24'd7655743, 24'd7710533, 24'd7899512, 24'd8185283, 24'd8511291, 24'd8813020, 24'd9030759, 24'd9121417, 24'd9067054, 24'd8878427, 24'd8592866, 24'd8266882, 24'd7964988, 24'd7746927, 24'd7655854, 24'd7709791, 24'd7898065, 24'd8183416, 24'd8509374, 24'd8811433, 
24'd9029815, 24'd9121304, 24'd9067793, 24'd8879873, 24'd8594732, 24'd8268800, 24'd7966577, 24'd7747873, 24'd7655970, 24'd7709054, 24'd7896621, 24'd8181551, 24'd8507457, 24'd8809843, 24'd9028867, 24'd9121185, 24'd9068528, 24'd8881315, 24'd8596597, 24'd8270717, 24'd7968169, 24'd7748824, 24'd7656091, 24'd7708322, 24'd7895180, 24'd8179687, 24'd8505538, 24'd8808250, 24'd9027914, 24'd9121062, 
24'd9069258, 24'd8882754, 24'd8598460, 24'd8272636, 24'd7969763, 24'd7749779, 24'd7656217, 24'd7707594, 24'd7893743, 24'd8177824, 24'd8503619, 24'd8806653, 24'd9026957, 24'd9120933, 24'd9069983, 24'd8884189, 24'd8600322, 24'd8274556, 24'd7971361, 24'd7750738, 24'd7656348, 24'd7706872, 24'd7892309, 24'd8175963, 24'd8501699, 24'd8805054, 24'd9025996, 24'd9120799, 24'd9070703, 24'd8885621, 
24'd8602182, 24'd8276476, 24'd7972961, 24'd7751702, 24'd7656485, 24'd7706154, 24'd7890879, 24'd8174104, 24'd8499778, 24'd8803453, 24'd9025030, 24'd9120660, 24'd9071418, 24'd8887050, 24'd8604040, 24'd8278397, 24'd7974565, 24'd7752670, 24'd7656627, 24'd7705441, 24'd7889452, 24'd8172246, 24'd8497857, 24'd8801848, 24'd9024059, 24'd9120516, 24'd9072129, 24'd8888475, 24'd8605898, 24'd8280319, 
24'd7976171, 24'd7753643, 24'd7656773, 24'd7704732, 24'd7888029, 24'd8170389, 24'd8495934, 24'd8800240, 24'd9023084, 24'd9120366, 24'd9072835, 24'd8889896, 24'd8607753, 24'd8282242, 24'd7977780, 24'd7754620, 24'd7656925, 24'd7704029, 24'd7886609, 24'd8168534, 24'd8494011, 24'd8798629, 24'd9022105, 24'd9120212, 24'd9073536, 24'd8891314, 24'd8609608, 24'd8284165, 24'd7979392, 24'd7755602, 
24'd7657082, 24'd7703330, 24'd7885193, 24'd8166681, 24'd8492088, 24'd8797016, 24'd9021121, 24'd9120052, 24'd9074233, 24'd8892729, 24'd8611460, 24'd8286090, 24'd7981007, 24'd7756588, 24'd7657244, 24'd7702636, 24'd7883780, 24'd8164829, 24'd8490163, 24'd8795399, 24'd9020132, 24'd9119888, 24'd9074924, 24'd8894140, 24'd8613311, 24'd8288014, 24'd7982625, 24'd7757578, 24'd7657412, 24'd7701947, 
24'd7882371, 24'd8162979, 24'd8488238, 24'd8793780, 24'd9019140, 24'd9119718, 24'd9075611, 24'd8895547, 24'd8615161, 24'd8289940, 24'd7984245, 24'd7758573, 24'd7657584, 24'd7701263, 24'd7880966, 24'd8161130, 24'd8486312, 24'd8792158, 24'd9018142, 24'd9119543, 24'd9076293, 24'd8896951, 24'd8617009, 24'd8291866, 24'd7985869, 24'd7759573, 24'd7657761, 24'd7700583, 24'd7879564, 24'd8159283, 
24'd8484385, 24'd8790533, 24'd9017141, 24'd9119363, 24'd9076970, 24'd8898351, 24'd8618855, 24'd8293793, 24'd7987495, 24'd7760577, 24'd7657944, 24'd7699909, 24'd7878165, 24'd8157438, 24'd8482458, 24'd8788906, 24'd9016135, 24'd9119178, 24'd9077642, 24'd8899748, 24'd8620700, 24'd8295721, 24'd7989124, 24'd7761585, 24'd7658132, 24'd7699239, 24'd7876770, 24'd8155594, 24'd8480530, 24'd8787275, 
24'd9015125, 24'd9118987, 24'd9078309, 24'd8901141, 24'd8622543, 24'd8297649, 24'd7990756, 24'd7762597, 24'd7658325, 24'd7698574, 24'd7875379, 24'd8153752, 24'd8478601, 24'd8785642, 24'd9014110, 24'd9118792, 24'd9078972, 24'd8902530, 24'd8624384, 24'd8299578, 24'd7992391, 24'd7763614, 24'd7658523, 24'd7697914, 24'd7873991, 24'd8151911, 24'd8476672, 24'd8784006, 24'd9013091, 24'd9118591, 
24'd9079630, 24'd8903916, 24'd8626224, 24'd8301508, 24'd7994028, 24'd7764636, 24'd7658726, 24'd7697258, 24'd7872607, 24'd8150072, 24'd8474742, 24'd8782367, 24'd9012067, 24'd9118386, 24'd9080283, 24'd8905298, 24'd8628062, 24'd8303438, 24'd7995669, 24'd7765661, 24'd7658934, 24'd7696608, 24'd7871227, 24'd8148235, 24'd8472812, 24'd8780725, 24'd9011039, 24'd9118175, 24'd9080931, 24'd8906677, 
24'd8629898, 24'd8305369, 24'd7997312, 24'd7766691, 24'd7659147, 24'd7695962, 24'd7869850, 24'd8146399, 24'd8470881, 24'd8779081, 24'd9010007, 24'd9117959, 24'd9081574, 24'd8908052, 24'd8631733, 24'd8307300, 24'd7998957, 24'd7767726, 24'd7659366, 24'd7695321, 24'd7868477, 24'd8144565, 24'd8468949, 24'd8777434, 24'd9008970, 24'd9117738, 24'd9082212, 24'd8909423, 24'd8633566, 24'd8309232, 
24'd8000606, 24'd7768765, 24'd7659589, 24'd7694685, 24'd7867107, 24'd8142733, 24'd8467017, 24'd8775784, 24'd9007929, 24'd9117512, 24'd9082846, 24'd8910791, 24'd8635397, 24'd8311164, 24'd8002257, 24'd7769808, 24'd7659818, 24'd7694054, 24'd7865741, 24'd8140903, 24'd8465084, 24'd8774131, 24'd9006884, 24'd9117281, 24'd9083474, 24'd8912155, 24'd8637227, 24'd8313097, 24'd8003911, 24'd7770855, 
24'd7660052, 24'd7693428, 24'd7864379, 24'd8139074, 24'd8463151, 24'd8772476, 24'd9005834, 24'd9117044, 24'd9084098, 24'd8913515, 24'd8639055, 24'd8315031, 24'd8005568, 24'd7771907, 24'd7660291, 24'd7692807, 24'd7863021, 24'd8137247, 24'd8461217, 24'd8770818, 24'd9004780, 24'd9116803, 24'd9084717, 24'd8914872, 24'd8640881, 24'd8316965, 24'd8007227, 24'd7772963, 24'd7660535, 24'd7692191, 
24'd7861666, 24'd8135422, 24'd8459283, 24'd8769158, 24'd9003722, 24'd9116556, 24'd9085331, 24'd8916225, 24'd8642705, 24'd8318899, 24'd8008889, 24'd7774024, 24'd7660784, 24'd7691579, 24'd7860315, 24'd8133599, 24'd8457348, 24'd8767494, 24'd9002659, 24'd9116305, 24'd9085940, 24'd8917574, 24'd8644527, 24'd8320834, 24'd8010553, 24'd7775089, 24'd7661038, 24'd7690972, 24'd7858967, 24'd8131777, 
24'd8455413, 24'd8765828, 24'd9001592, 24'd9116048, 24'd9086544, 24'd8918920, 24'd8646348, 24'd8322770, 24'd8012221, 24'd7776158, 24'd7661298, 24'd7690371, 24'd7857623, 24'd8129957, 24'd8453477, 24'd8764160, 24'd9000521, 24'd9115786, 24'd9087143, 24'd8920262, 24'd8648167, 24'd8324706, 24'd8013891, 24'd7777231, 24'd7661562, 24'd7689774, 24'd7856283, 24'd8128139, 24'd8451541, 24'd8762488, 
24'd8999446, 24'd9115519, 24'd9087738, 24'd8921600, 24'd8649984, 24'd8326642, 24'd8015563, 24'd7778309, 24'd7661831, 24'd7689182, 24'd7854947, 24'd8126323, 24'd8449604, 24'd8760815, 24'd8998366, 24'd9115247, 24'd9088327, 24'd8922935, 24'd8651799, 24'd8328579, 24'd8017238, 24'd7779391, 24'd7662106, 24'd7688595, 24'd7853615, 24'd8124509, 24'd8447667, 24'd8759138, 24'd8997282, 24'd9114970, 
24'd9088912, 24'd8924265, 24'd8653613, 24'd8330516, 24'd8018916, 24'd7780477, 24'd7662386, 24'd7688013, 24'd7852286, 24'd8122696, 24'd8445730, 24'd8757459, 24'd8996193, 24'd9114687, 24'd9089492, 24'd8925592, 24'd8655424, 24'd8332454, 24'd8020596, 24'd7781567, 24'd7662671, 24'd7687435, 24'd7850961, 24'd8120886, 24'd8443792, 24'd8755777, 24'd8995101, 24'd9114400, 24'd9090066, 24'd8926915, 
24'd8657234, 24'd8334392, 24'd8022279, 24'd7782662, 24'd7662960, 24'd7686863, 24'd7849640, 24'd8119077, 24'd8441854, 24'd8754093, 24'd8994004, 24'd9114108, 24'd9090636, 24'd8928235, 24'd8659042, 24'd8336331, 24'd8023965, 24'd7783761, 24'd7663255, 24'd7686296, 24'd7848322, 24'd8117270, 24'd8439915, 24'd8752406, 24'd8992903, 24'd9113810, 24'd9091201, 24'd8929550, 24'd8660848, 24'd8338269, 
24'd8025653, 24'd7784864, 24'd7663556, 24'd7685733, 24'd7847008, 24'd8115465, 24'd8437976, 24'd8750717, 24'd8991797, 24'd9113508, 24'd9091761, 24'd8930862, 24'd8662652, 24'd8340209, 24'd8027343, 24'd7785972, 24'd7663861, 24'd7685176, 24'd7845698, 24'd8113662, 24'd8436037, 24'd8749025, 24'd8990688, 24'd9113200, 24'd9092316, 24'd8932170, 24'd8664454, 24'd8342148, 24'd8029037, 24'd7787084, 
24'd7664171, 24'd7684623, 24'd7844392, 24'd8111861, 24'd8434097, 24'd8747331, 24'd8989574, 24'd9112887, 24'd9092866, 24'd8933474, 24'd8666254, 24'd8344088, 24'd8030732, 24'd7788199, 24'd7664486, 24'd7684075, 24'd7843090, 24'd8110062, 24'd8432157, 24'd8745634, 24'd8988456, 24'd9112569, 24'd9093412, 24'd8934775, 24'd8668052, 24'd8346028, 24'd8032430, 24'd7789320, 24'd7664807, 24'd7683533, 
24'd7841792, 24'd8108264, 24'd8430217, 24'd8743935, 24'd8987334, 24'd9112246, 24'd9093952, 24'd8936071, 24'd8669848, 24'd8347969, 24'd8034131, 24'd7790444, 24'd7665132, 24'd7682995, 24'd7840497, 24'd8106469, 24'd8428276, 24'd8742233, 24'd8986207, 24'd9111918, 24'd9094487, 24'd8937364, 24'd8671643, 24'd8349909, 24'd8035834, 24'd7791572, 24'd7665463, 24'd7682462, 24'd7839206, 24'd8104676, 
24'd8426335, 24'd8740528, 24'd8985077, 24'd9111585, 24'd9095018, 24'd8938653, 24'd8673435, 24'd8351850, 24'd8037540, 24'd7792705, 24'd7665798, 24'd7681934, 24'd7837919, 24'd8102885, 24'd8424394, 24'd8738821, 24'd8983942, 24'd9111247, 24'd9095543, 24'd8939938, 24'd8675225, 24'd8353792, 24'd8039248, 24'd7793842, 24'd7666139, 24'd7681411, 24'd7836636, 24'd8101095, 24'd8422453, 24'd8737112, 
24'd8982803, 24'd9110904, 24'd9096063, 24'd8941219, 24'd8677013, 24'd8355733, 24'd8040958, 24'd7794983, 24'd7666485, 24'd7680893, 24'd7835357, 24'd8099308, 24'd8420511, 24'd8735400, 24'd8981660, 24'd9110556, 24'd9096579, 24'd8942496, 24'd8678800, 24'd8357675, 24'd8042671, 24'd7796128, 24'd7666835, 24'd7680380, 24'd7834082, 24'd8097523, 24'd8418569, 24'd8733686, 24'd8980513, 24'd9110202, 
24'd9097090, 24'd8943770, 24'd8680584, 24'd8359617, 24'd8044387, 24'd7797277, 24'd7667191, 24'd7679872, 24'd7832810, 24'd8095740, 24'd8416627, 24'd8731970, 24'd8979361, 24'd9109844, 24'd9097595, 24'd8945039, 24'd8682366, 24'd8361559, 24'd8046105, 24'd7798431, 24'd7667552, 24'd7679369, 24'd7831543, 24'd8093959, 24'd8414685, 24'd8730251, 24'd8978206, 24'd9109480, 24'd9098096, 24'd8946305, 
24'd8684146, 24'd8363501, 24'd8047825, 24'd7799589, 24'd7667918, 24'd7678871, 24'd7830279, 24'd8092180, 24'd8412742, 24'd8728529, 24'd8977046, 24'd9109112, 24'd9098591, 24'd8947566, 24'd8685924, 24'd8365444, 24'd8049547, 24'd7800750, 24'd7668289, 24'd7678378, 24'd7829019, 24'd8090403, 24'd8410800, 24'd8726805, 24'd8975882, 24'd9108738, 24'd9099082, 24'd8948824, 24'd8687700, 24'd8367386, 
24'd8051272, 24'd7801916, 24'd7668665, 24'd7677890, 24'd7827764, 24'd8088628, 24'd8408857, 24'd8725079, 24'd8974714, 24'd9108360, 24'd9099568, 24'd8950078, 24'd8689474, 24'd8369329, 24'd8053000, 24'd7803086, 24'd7669046, 24'd7677406, 24'd7826512, 24'd8086855, 24'd8406914, 24'd8723351, 24'd8973542, 24'd9107976, 24'd9100048, 24'd8951328, 24'd8691246, 24'd8371272, 24'd8054729, 24'd7804260, 
24'd7669433, 24'd7676928, 24'd7825264, 24'd8085084, 24'd8404971, 24'd8721620, 24'd8972366, 24'd9107587, 24'd9100524, 24'd8952574, 24'd8693015, 24'd8373215, 24'd8056461, 24'd7805439, 24'd7669824, 24'd7676455, 24'd7824020, 24'd8083316, 24'd8403028, 24'd8719887, 24'd8971186, 24'd9107194, 24'd9100995, 24'd8953816, 24'd8694783, 24'd8375159, 24'd8058196, 24'd7806621, 24'd7670220, 24'd7675987, 
24'd7822780, 24'd8081549, 24'd8401085, 24'd8718151, 24'd8970001, 24'd9106795, 24'd9101460, 24'd8955054, 24'd8696548, 24'd8377102, 24'd8059933, 24'd7807807, 24'd7670621, 24'd7675524, 24'd7821544, 24'd8079785, 24'd8399141, 24'd8716413, 24'd8968813, 24'd9106391, 24'd9101921, 24'd8956288, 24'd8698311, 24'd8379045, 24'd8061671, 24'd7808998, 24'd7671028, 24'd7675065, 24'd7820312, 24'd8078023, 
24'd8397198, 24'd8714673, 24'd8967621, 24'd9105982, 24'd9102377, 24'd8957518, 24'd8700072, 24'd8380989, 24'd8063413, 24'd7810192, 24'd7671439, 24'd7674612, 24'd7819084, 24'd8076263, 24'd8395255, 24'd8712931, 24'd8966424, 24'd9105568, 24'd9102828, 24'd8958744, 24'd8701831, 24'd8382932, 24'd8065156, 24'd7811391, 24'd7671855, 24'd7674164, 24'd7817860, 24'd8074505, 24'd8393311, 24'd8711186, 
24'd8965223, 24'd9105149, 24'd9103273, 24'd8959966, 24'd8703588, 24'd8384876, 24'd8066902, 24'd7812593, 24'd7672277, 24'd7673721, 24'd7816640, 24'd8072750, 24'd8391367, 24'd8709439, 24'd8964019, 24'd9104726, 24'd9103714, 24'd8961184, 24'd8705342, 24'd8386819, 24'd8068650, 24'd7813800, 24'd7672703, 24'd7673283, 24'd7815423, 24'd8070996, 24'd8389424, 24'd8707690, 24'd8962810, 24'd9104297, 
24'd9104150, 24'd8962398, 24'd8707094, 24'd8388763, 24'd8070401, 24'd7815011, 24'd7673135, 24'd7672849, 24'd7814211, 24'd8069245, 24'd8387480, 24'd8705938, 24'd8961597, 24'd9103863, 24'd9104580, 24'd8963608, 24'd8708844, 24'd8390706, 24'd8072153, 24'd7816225, 24'd7673571, 24'd7672421, 24'd7813003, 24'd8067496, 24'd8385537, 24'd8704185, 24'd8960381, 24'd9103424, 24'd9105006, 24'd8964814, 
24'd8710592, 24'd8392650, 24'd8073908, 24'd7817444, 24'd7674013, 24'd7671998, 24'd7811799, 24'd8065750, 24'd8383593, 24'd8702429, 24'd8959160, 24'd9102980, 24'd9105426, 24'd8966016, 24'd8712338, 24'd8394594, 24'd8075665, 24'd7818667, 24'd7674459, 24'd7671580, 24'd7810599, 24'd8064005, 24'd8381650, 24'd8700671, 24'd8957935, 24'd9102531, 24'd9105842, 24'd8967214, 24'd8714081, 24'd8396537, 
24'd8077424, 24'd7819894, 24'd7674911, 24'd7671167, 24'd7809404, 24'd8062263, 24'd8379706, 24'd8698911, 24'd8956706, 24'd9102077, 24'd9106253, 24'd8968408, 24'd8715822, 24'd8398480, 24'd8079185, 24'd7821124, 24'd7675367, 24'd7670759, 24'd7808212, 24'd8060524, 24'd8377763, 24'd8697148, 24'd8955474, 24'd9101618, 24'd9106658, 24'd8969598, 24'd8717560, 24'd8400424, 24'd8080949, 24'd7822359, 
24'd7675829, 24'd7670356, 24'd7807024, 24'd8058786, 24'd8375820, 24'd8695384, 24'd8954237, 24'd9101154, 24'd9107059, 24'd8970783, 24'd8719297, 24'd8402367, 24'd8082715, 24'd7823598, 24'd7676295, 24'd7669958, 24'd7805840, 24'd8057051, 24'd8373876, 24'd8693617, 24'd8952996, 24'd9100685, 24'd9107454, 24'd8971965, 24'd8721031, 24'd8404310, 24'd8084482, 24'd7824840, 24'd7676767, 24'd7669565, 
24'd7804661, 24'd8055318, 24'd8371933, 24'd8691848, 24'd8951752, 24'd9100211, 24'd9107844, 24'd8973143, 24'd8722762, 24'd8406253, 24'd8086252, 24'd7826087, 24'd7677243, 24'd7669177, 24'd7803485, 24'd8053588, 24'd8369990, 24'd8690077, 24'd8950503, 24'd9099732, 24'd9108230, 24'd8974316, 24'd8724492, 24'd8408196, 24'd8088024, 24'd7827337, 24'd7677725, 24'd7668794, 24'd7802314, 24'd8051860, 
24'd8368047, 24'd8688304, 24'd8949251, 24'd9099248, 24'd9108610, 24'd8975485, 24'd8726219, 24'd8410139, 24'd8089799, 24'd7828592, 24'd7678211, 24'd7668417, 24'd7801146, 24'd8050134, 24'd8366104, 24'd8686528, 24'd8947994, 24'd9098759, 24'd9108985, 24'd8976651, 24'd8727943, 24'd8412082, 24'd8091575, 24'd7829850, 24'd7678703, 24'd7668044, 24'd7799983, 24'd8048410, 24'd8364162, 24'd8684751, 
24'd8946734, 24'd9098265, 24'd9109356, 24'd8977812, 24'd8729665, 24'd8414024, 24'd8093353, 24'd7831113, 24'd7679199, 24'd7667676, 24'd7798824, 24'd8046689, 24'd8362219, 24'd8682972, 24'd8945470, 24'd9097766, 24'd9109721, 24'd8978969, 24'd8731385, 24'd8415967, 24'd8095134, 24'd7832379, 24'd7679700, 24'd7667313, 24'd7797669, 24'd8044971, 24'd8360277, 24'd8681190, 24'd8944202, 24'd9097262, 
24'd9110081, 24'd8980122, 24'd8733103, 24'd8417909, 24'd8096916, 24'd7833649, 24'd7680207, 24'd7666956, 24'd7796519, 24'd8043255, 24'd8358335, 24'd8679407, 24'd8942930, 24'd9096753, 24'd9110436, 24'd8981270, 24'd8734818, 24'd8419851, 24'd8098701, 24'd7834923, 24'd7680718, 24'd7666603, 24'd7795372, 24'd8041541, 24'd8356393, 24'd8677621, 24'd8941654, 24'd9096239, 24'd9110786, 24'd8982415, 
24'd8736530, 24'd8421792, 24'd8100487, 24'd7836201, 24'd7681234, 24'd7666256, 24'd7794230, 24'd8039829, 24'd8354452, 24'd8675834, 24'd8940374, 24'd9095721, 24'd9111131, 24'd8983555, 24'd8738240, 24'd8423734, 24'd8102276, 24'd7837482, 24'd7681756, 24'd7665914, 24'd7793091, 24'd8038120, 24'd8352510, 24'd8674044, 24'd8939090, 24'd9095197, 24'd9111471, 24'd8984691, 24'd8739948, 24'd8425675, 
24'd8104067, 24'd7838768, 24'd7682282, 24'd7665576, 24'd7791957, 24'd8036414, 24'd8350569, 24'd8672252, 24'd8937803, 24'd9094668, 24'd9111806, 24'd8985823, 24'd8741653, 24'd8427616, 24'd8105859, 24'd7840058, 24'd7682813, 24'd7665244, 24'd7790827, 24'd8034710, 24'd8348629, 24'd8670459, 24'd8936511, 24'd9094135, 24'd9112135, 24'd8986951, 24'd8743356, 24'd8429557, 24'd8107654, 24'd7841351, 
24'd7683349, 24'd7664917, 24'd7789701, 24'd8033009, 24'd8346688, 24'd8668663, 24'd8935216, 24'd9093596, 24'd9112460, 24'd8988075, 24'd8745056, 24'd8431497, 24'd8109450, 24'd7842648, 24'd7683890, 24'd7664595, 24'd7788580, 24'd8031310, 24'd8344748, 24'd8666866, 24'd8933917, 24'd9093052, 24'd9112780, 24'd8989194, 24'd8746754, 24'd8433437, 24'd8111249, 24'd7843949, 24'd7684436, 24'd7664278, 
24'd7787463, 24'd8029613, 24'd8342808, 24'd8665066, 24'd8932614, 24'd9092504, 24'd9113094, 24'd8990310, 24'd8748449, 24'd8435377, 24'd8113049, 24'd7845254, 24'd7684987, 24'd7663966, 24'd7786349, 24'd8027919, 24'd8340868, 24'd8663265, 24'd8931307, 24'd9091951, 24'd9113403, 24'd8991421, 24'd8750142, 24'd8437317, 24'd8114852, 24'd7846562, 24'd7685543, 24'd7663659, 24'd7785241, 24'd8026228, 
24'd8338929, 24'd8661462, 24'd8929997, 24'd9091392, 24'd9113708, 24'd8992527, 24'd8751832, 24'd8439256, 24'd8116656, 24'd7847875, 24'd7686104, 24'd7663357, 24'd7784136, 24'd8024539, 24'd8336990, 24'd8659656, 24'd8928683, 24'd9090829, 24'd9114007, 24'd8993630, 24'd8753520, 24'd8441194, 24'd8118462, 24'd7849191, 24'd7686670, 24'd7663060, 24'd7783035, 24'd8022852, 24'd8335051, 24'd8657849, 
24'd8927364, 24'd9090261, 24'd9114301, 24'd8994728, 24'd8755205, 24'd8443133, 24'd8120270, 24'd7850511, 24'd7687240, 24'd7662769, 24'd7781939, 24'd8021168, 24'd8333113, 24'd8656040, 24'd8926043, 24'd9089688, 24'd9114590, 24'd8995822, 24'd8756887, 24'd8445071, 24'd8122080, 24'd7851835, 24'd7687816, 24'd7662482, 24'd7780847, 24'd8019487, 24'd8331175, 24'd8654229, 24'd8924717, 24'd9089110, 
24'd9114874, 24'd8996912, 24'd8758567, 24'd8447008, 24'd8123892, 24'd7853162, 24'd7688396, 24'd7662201, 24'd7779760, 24'd8017809, 24'd8329238, 24'd8652416, 24'd8923388, 24'd9088527, 24'd9115153, 24'd8997998, 24'd8760245, 24'd8448946, 24'd8125706, 24'd7854494, 24'd7688982, 24'd7661924, 24'd7778676, 24'd8016133, 24'd8327301, 24'd8650602, 24'd8922054, 24'd9087939, 24'd9115427, 24'd8999079, 
24'd8761919, 24'd8450882, 24'd8127521, 24'd7855829, 24'd7689572, 24'd7661653, 24'd7777597, 24'd8014459, 24'd8325364, 24'd8648785, 24'd8920718, 24'd9087346, 24'd9115696, 24'd9000156, 24'd8763592, 24'd8452819, 24'd8129339, 24'd7857167, 24'd7690167, 24'd7661387, 24'd7776522, 24'd8012788, 24'd8323428, 24'd8646967, 24'd8919377, 24'd9086748, 24'd9115959, 24'd9001228, 24'd8765261, 24'd8454755, 
24'd8131158, 24'd7858510, 24'd7690767, 24'd7661126, 24'd7775452, 24'd8011120, 24'd8321493, 24'd8645147, 24'd8918033, 24'd9086146, 24'd9116218, 24'd9002297, 24'd8766928, 24'd8456690, 24'd8132979, 24'd7859856, 24'd7691372, 24'd7660870, 24'd7774386, 24'd8009455, 24'd8319557, 24'd8643325, 24'd8916684, 24'd9085539, 24'd9116471, 24'd9003361, 24'd8768592, 24'd8458625, 24'd8134802, 24'd7861206, 
24'd7691982, 24'd7660619, 24'd7773324, 24'd8007792, 24'd8317623, 24'd8641501, 24'd8915333, 24'd9084926, 24'd9116720, 24'd9004421, 24'd8770254, 24'd8460560, 24'd8136626, 24'd7862560, 24'd7692597, 24'd7660373, 24'd7772266, 24'd8006132, 24'd8315688, 24'd8639676, 24'd8913977, 24'd9084309, 24'd9116963, 24'd9005476, 24'd8771913, 24'd8462493, 24'd8138453, 24'd7863917, 24'd7693216, 24'd7660133, 
24'd7771213, 24'd8004474, 24'd8313755, 24'd8637849, 24'd8912618, 24'd9083687, 24'd9117201, 24'd9006527, 24'd8773569, 24'd8464427, 24'd8140281, 24'd7865278, 24'd7693841, 24'd7659897, 24'd7770164, 24'd8002819, 24'd8311822, 24'd8636020, 24'd8911255, 24'd9083060, 24'd9117434, 24'd9007574, 24'd8775222, 24'd8466360, 24'd8142110, 24'd7866642, 24'd7694470, 24'd7659667, 24'd7769119, 24'd8001167, 
24'd8309889, 24'd8634189, 24'd8909889, 24'd9082428, 24'd9117662, 24'd9008617, 24'd8776873, 24'd8468292, 24'd8143942, 24'd7868011, 24'd7695105, 24'd7659441, 24'd7768079, 24'd7999518, 24'd8307957, 24'd8632357, 24'd8908519, 24'd9081792, 24'd9117884, 24'd9009655, 24'd8778521, 24'd8470224, 24'd8145775, 24'd7869383, 24'd7695744, 24'd7659221, 24'd7767043, 24'd7997871, 24'd8306025, 24'd8630522, 
24'd8907145, 24'd9081150, 24'd9118102, 24'd9010689, 24'd8780166, 24'd8472155, 24'd8147610, 24'd7870758, 24'd7696388, 24'd7659006, 24'd7766011, 24'd7996227, 24'd8304094, 24'd8628687, 24'd8905768, 24'd9080504, 24'd9118315, 24'd9011718, 24'd8781809, 24'd8474086, 24'd8149447, 24'd7872137, 24'd7697036, 24'd7658796, 24'd7764984, 24'd7994586, 24'd8302164, 24'd8626849, 24'd8904387, 24'd9079852, 
24'd9118522, 24'd9012743, 24'd8783449, 24'd8476016, 24'd8151285, 24'd7873520, 24'd7697690, 24'd7658591, 24'd7763961, 24'd7992948, 24'd8300234, 24'd8625010, 24'd8903002, 24'd9079196, 24'd9118724, 24'd9013764, 24'd8785086, 24'd8477945, 24'd8153125, 24'd7874907, 24'd7698349, 24'd7658391, 24'd7762943, 24'd7991312, 24'd8298305, 24'd8623169, 24'd8901614, 24'd9078535, 24'd9118921, 24'd9014780, 
24'd8786720, 24'd8479874, 24'd8154967, 24'd7876297, 24'd7699012, 24'd7658197, 24'd7761929, 24'd7989679, 24'd8296377, 24'd8621327, 24'd8900222, 24'd9077870, 24'd9119114, 24'd9015792, 24'd8788351, 24'd8481802, 24'd8156810, 24'd7877690, 24'd7699680, 24'd7658007, 24'd7760919, 24'd7988049, 24'd8294449, 24'd8619482, 24'd8898826, 24'd9077199, 24'd9119300, 24'd9016799, 24'd8789980, 24'd8483730, 
24'd8158655, 24'd7879088, 24'd7700353, 24'd7657823, 24'd7759914, 24'd7986422, 24'd8292522, 24'd8617637, 24'd8897427, 24'd9076523, 24'd9119482, 24'd9017802, 24'd8791606, 24'd8485657, 24'd8160502, 24'd7880489, 24'd7701031, 24'd7657644, 24'd7758913, 24'd7984797, 24'd8290595, 24'd8615789, 24'd8896025, 24'd9075843, 24'd9119659, 24'd9018801, 24'd8793229, 24'd8487583, 24'd8162350, 24'd7881893, 
24'd7701714, 24'd7657470, 24'd7757916, 24'd7983176, 24'd8288669, 24'd8613940, 24'd8894619, 24'd9075158, 24'd9119831, 24'd9019795, 24'd8794849, 24'd8489508, 24'd8164200, 24'd7883301, 24'd7702401, 24'd7657301, 24'd7756924, 24'd7981557, 24'd8286744, 24'd8612090, 24'd8893209, 24'd9074468, 24'd9119997, 24'd9020785, 24'd8796466, 24'd8491433, 24'd8166051, 24'd7884712, 24'd7703093, 24'd7657137, 
24'd7755937, 24'd7979941, 24'd8284820, 24'd8610238, 24'd8891796, 24'd9073774, 24'd9120158, 24'd9021770, 24'd8798081, 24'd8493357, 24'd8167904, 24'd7886127, 24'd7703791, 24'd7656978, 24'd7754953, 24'd7978328, 24'd8282896, 24'd8608384, 24'd8890379, 24'd9073074, 24'd9120314, 24'd9022751, 24'd8799692, 24'd8495281, 24'd8169758, 24'd7887546, 24'd7704492, 24'd7656824, 24'd7753975, 24'd7976718, 
24'd8280973, 24'd8606529, 24'd8888959, 24'd9072370, 24'd9120466, 24'd9023728, 24'd8801301, 24'd8497203, 24'd8171614, 24'd7888968, 24'd7705199, 24'd7656676, 24'd7753000, 24'd7975111, 24'd8279051, 24'd8604672, 24'd8887535, 24'd9071661, 24'd9120611, 24'd9024700, 24'd8802907, 24'd8499125, 24'd8173472, 24'd7890393, 24'd7705911, 24'd7656533, 24'd7752031, 24'd7973506, 24'd8277129, 24'd8602814, 
24'd8886108, 24'd9070947, 24'd9120752, 24'd9025668, 24'd8804510, 24'd8501046, 24'd8175331, 24'd7891822, 24'd7706627, 24'd7656394, 24'd7751065, 24'd7971905, 24'd8275209, 24'd8600954, 24'd8884677, 24'd9070228, 24'd9120888, 24'd9026631, 24'd8806110, 24'd8502966, 24'd8177191, 24'd7893255, 24'd7707348, 24'd7656261, 24'd7750104, 24'd7970306, 24'd8273289, 24'd8599093, 24'd8883243, 24'd9069505, 
24'd9121018, 24'd9027589, 24'd8807707, 24'd8504886, 24'd8179053, 24'd7894691, 24'd7708074, 24'd7656133, 24'd7749148, 24'd7968711, 24'd8271370, 24'd8597230, 24'd8881805, 24'd9068776, 24'd9121144, 24'd9028544, 24'd8809301, 24'd8506804, 24'd8180916, 24'd7896130, 24'd7708804, 24'd7656010, 24'd7748196, 24'd7967118, 24'd8269452, 24'd8595366, 24'd8880364, 24'd9068043, 24'd9121264, 24'd9029493, 
24'd8810892, 24'd8508722, 24'd8182781, 24'd7897573, 24'd7709540, 24'd7655893, 24'd7747249, 24'd7965528, 24'd8267534, 24'd8593501, 24'd8878919, 24'd9067306, 24'd9121379, 24'd9030438, 24'd8812481, 24'd8510639, 24'd8184648, 24'd7899020, 24'd7710280, 24'd7655780, 24'd7746306, 24'd7963941, 24'd8265618, 24'd8591634, 24'd8877471, 24'd9066563, 24'd9121489, 24'd9031379, 24'd8814066, 24'd8512555, 
24'd8186515, 24'd7900469, 24'd7711025, 24'd7655673, 24'd7745367, 24'd7962358, 24'd8263702, 24'd8589765, 24'd8876020, 24'd9065816, 24'd9121594, 24'd9032315, 24'd8815648, 24'd8514470, 24'd8188385, 24'd7901922, 24'd7711775, 24'd7655571, 24'd7744433, 24'd7960777, 24'd8261787, 24'd8587895, 24'd8874565, 24'd9065064, 24'd9121694, 24'd9033247, 24'd8817227, 24'd8516385, 24'd8190255, 24'd7903379, 
24'd7712529, 24'd7655473, 24'd7743504, 24'd7959199, 24'd8259873, 24'd8586024, 24'd8873106, 24'd9064307, 24'd9121788, 24'd9034174, 24'd8818804, 24'd8518298, 24'd8192127, 24'd7904839, 24'd7713288, 24'd7655381, 24'd7742579, 24'd7957624, 24'd8257960, 24'd8584151, 24'd8871645, 24'd9063546, 24'd9121878, 24'd9035097, 24'd8820377, 24'd8520211, 24'd8194000, 24'd7906303, 24'd7714052, 24'd7655295, 
24'd7741659, 24'd7956053, 24'd8256048, 24'd8582277, 24'd8870180, 24'd9062779, 24'd9121962, 24'd9036015, 24'd8821947, 24'd8522122, 24'd8195875, 24'd7907769, 24'd7714820, 24'd7655213, 24'd7740743, 24'd7954484, 24'd8254137, 24'd8580402, 24'd8868711, 24'd9062008, 24'd9122041, 24'd9036928, 24'd8823514, 24'd8524033, 24'd8197751, 24'd7909239, 24'd7715594, 24'd7655136, 24'd7739831, 24'd7952918, 
24'd8252227, 24'd8578525, 24'd8867239, 24'd9061233, 24'd9122115, 24'd9037837, 24'd8825078, 24'd8525943, 24'd8199629, 24'd7910713, 24'd7716372, 24'd7655065, 24'd7738925, 24'd7951356, 24'd8250318, 24'd8576647, 24'd8865764, 24'd9060452, 24'd9122184, 24'd9038742, 24'd8826640, 24'd8527851, 24'd8201507, 24'd7912190, 24'd7717155, 24'd7654999, 24'd7738023, 24'd7949796, 24'd8248410, 24'd8574768, 
24'd8864285, 24'd9059667, 24'd9122248, 24'd9039642, 24'd8828198, 24'd8529759, 24'd8203387, 24'd7913670, 24'd7717942, 24'd7654938, 24'd7737125, 24'd7948240, 24'd8246502, 24'd8572887, 24'd8862804, 24'd9058877, 24'd9122306, 24'd9040537, 24'd8829753, 24'd8531666, 24'd8205269, 24'd7915154, 24'd7718734, 24'd7654882, 24'd7736232, 24'd7946686, 24'd8244596, 24'd8571005, 24'd8861318, 24'd9058083, 
24'd9122360, 24'd9041428, 24'd8831304, 24'd8533572, 24'd8207151, 24'd7916640, 24'd7719531, 24'd7654831, 24'd7735343, 24'd7945136, 24'd8242691, 24'd8569122, 24'd8859830, 24'd9057284, 24'd9122408, 24'd9042314, 24'd8832853, 24'd8535477, 24'd8209035, 24'd7918131, 24'd7720333, 24'd7654785, 24'd7734460, 24'd7943589, 24'd8240786, 24'd8567237, 24'd8858338, 24'd9056480, 24'd9122451, 24'd9043196, 
24'd8834399, 24'd8537380, 24'd8210920, 24'd7919624, 24'd7721139, 24'd7654744, 24'd7733580, 24'd7942045, 24'd8238883, 24'd8565352, 24'd8856843, 24'd9055671, 24'd9122489, 24'd9044073, 24'd8835941, 24'd8539283, 24'd8212807, 24'd7921121, 24'd7721950, 24'd7654709, 24'd7732705, 24'd7940504, 24'd8236981, 24'd8563465, 24'd8855345, 24'd9054858, 24'd9122522, 24'd9044945, 24'd8837481, 24'd8541185, 
24'd8214694, 24'd7922621, 24'd7722765, 24'd7654679, 24'd7731835, 24'd7938966, 24'd8235080, 24'd8561576, 24'd8853843, 24'd9054040, 24'd9122549, 24'd9045813, 24'd8839017, 24'd8543085, 24'd8216583, 24'd7924124, 24'd7723586, 24'd7654654, 24'd7730970, 24'd7937431, 24'd8233180, 24'd8559687, 24'd8852338, 24'd9053218, 24'd9122572, 24'd9046676, 24'd8840550, 24'd8544985, 24'd8218473, 24'd7925631, 
24'd7724411, 24'd7654634, 24'd7730109, 24'd7935900, 24'd8231281, 24'd8557796, 24'd8850830, 24'd9052390, 24'd9122589, 24'd9047535, 24'd8842080, 24'd8546883, 24'd8220364, 24'd7927141, 24'd7725240, 24'd7654619, 24'd7729253, 24'd7934372, 24'd8229383, 24'd8555905, 24'd8849318, 24'd9051558, 24'd9122602, 24'd9048389, 24'd8843606, 24'd8548781, 24'd8222257, 24'd7928654, 24'd7726074, 24'd7654609, 
24'd7728401, 24'd7932846, 24'd8227486, 24'd8554012, 24'd8847804, 24'd9050722, 24'd9122609, 24'd9049238, 24'd8845130, 24'd8550677, 24'd8224150, 24'd7930170, 24'd7726913, 24'd7654605, 24'd7727554, 24'd7931325, 24'd8225591, 24'd8552117, 24'd8846286, 24'd9049881, 24'd9122611, 24'd9050083, 24'd8846650, 24'd8552572, 24'd8226045, 24'd7931689, 24'd7727757, 24'd7654605, 24'd7726712, 24'd7929806, 
24'd8223696, 24'd8550222, 24'd8844765, 24'd9049035, 24'd9122607, 24'd9050923, 24'd8848167, 24'd8554466, 24'd8227941, 24'd7933212, 24'd7728605, 24'd7654611, 24'd7725874, 24'd7928290, 24'd8221803, 24'd8548326, 24'd8843240, 24'd9048184, 24'd9122599, 24'd9051758, 24'd8849681, 24'd8556358, 24'd8229838, 24'd7934738, 24'd7729458, 24'd7654622, 24'd7725041, 24'd7926778, 24'd8219911, 24'd8546428, 
24'd8841713, 24'd9047329, 24'd9122586, 24'd9052589, 24'd8851192, 24'd8558250, 24'd8231736, 24'd7936267, 24'd7730315, 24'd7654638, 24'd7724212, 24'd7925269, 24'd8218020, 24'd8544529, 24'd8840182, 24'd9046470, 24'd9122567, 24'd9053415, 24'd8852699, 24'd8560140, 24'd8233635, 24'd7937799, 24'd7731177, 24'd7654659, 24'd7723388, 24'd7923763, 24'd8216130, 24'd8542630, 24'd8838649, 24'd9045605, 
24'd9122543, 24'd9054237, 24'd8854203, 24'd8562029, 24'd8235536, 24'd7939335, 24'd7732044, 24'd7654686, 24'd7722569, 24'd7922261, 24'd8214241, 24'd8540729, 24'd8837112, 24'd9044736, 24'd9122514, 24'd9055054, 24'd8855704, 24'd8563917, 24'd8237437, 24'd7940873, 24'd7732915, 24'd7654717, 24'd7721755, 24'd7920762, 24'd8212354, 24'd8538827, 24'd8835572, 24'd9043863, 24'd9122480, 24'd9055866, 
24'd8857202, 24'd8565804, 24'd8239339, 24'd7942415, 24'd7733791, 24'd7654754, 24'd7720945, 24'd7919266, 24'd8210468, 24'd8536924, 24'd8834028, 24'd9042985, 24'd9122441, 24'd9056673, 24'd8858696, 24'd8567690, 24'd8241243, 24'd7943960, 24'd7734671, 24'd7654795, 24'd7720140, 24'd7917773, 24'd8208583, 24'd8535020, 24'd8832482, 24'd9042102, 24'd9122397, 24'd9057476, 24'd8860187, 24'd8569574, 
24'd8243147, 24'd7945507, 24'd7735556, 24'd7654842, 24'd7719340, 24'd7916284, 24'd8206700, 24'd8533115, 24'd8830932, 24'd9041215, 24'd9122347, 24'd9058274, 24'd8861675, 24'd8571457, 24'd8245053, 24'd7947058, 24'd7736446, 24'd7654894, 24'd7718544, 24'd7914797, 24'd8204817, 24'd8531209, 24'd8829380, 24'd9040323, 24'd9122293, 24'd9059067, 24'd8863159, 24'd8573338, 24'd8246960, 24'd7948613, 
24'd7737340, 24'd7654952, 24'd7717753, 24'd7913315, 24'd8202936, 24'd8529302, 24'd8827824, 24'd9039426, 24'd9122233, 24'd9059856, 24'd8864640, 24'd8575219, 24'd8248867, 24'd7950170, 24'd7738239, 24'd7655014, 24'd7716966, 24'd7911835, 24'd8201057, 24'd8527394, 24'd8826265, 24'd9038525, 24'd9122168, 24'd9060640, 24'd8866118, 24'd8577098, 24'd8250776, 24'd7951730, 24'd7739142, 24'd7655082, 
24'd7716185, 24'd7910359, 24'd8199178, 24'd8525485, 24'd8824704, 24'd9037620, 24'd9122098, 24'd9061419, 24'd8867593, 24'd8578976, 24'd8252685, 24'd7953293, 24'd7740050, 24'd7655154, 24'd7715408, 24'd7908887, 24'd8197301, 24'd8523575, 24'd8823139, 24'd9036710, 24'd9122023, 24'd9062194, 24'd8869064, 24'd8580852, 24'd8254596, 24'd7954860, 24'd7740962, 24'd7655232, 24'd7714636, 24'd7907417, 
24'd8195425, 24'd8521664, 24'd8821571, 24'd9035795, 24'd9121942, 24'd9062964, 24'd8870531, 24'd8582727, 24'd8256507, 24'd7956429, 24'd7741879, 24'd7655315, 24'd7713868, 24'd7905951, 24'd8193551, 24'd8519752, 24'd8820000, 24'd9034876, 24'd9121857, 24'd9063729, 24'd8871996, 24'd8584601, 24'd8258419, 24'd7958002, 24'd7742800, 24'd7655403, 24'd7713106, 24'd7904489, 24'd8191678, 24'd8517839, 
24'd8818426, 24'd9033952, 24'd9121766, 24'd9064489, 24'd8873456, 24'd8586473, 24'd8260332, 24'd7959577, 24'd7743726, 24'd7655496, 24'd7712348, 24'd7903029, 24'd8189806, 24'd8515926, 24'd8816849, 24'd9033024, 24'd9121670, 24'd9065245, 24'd8874914, 24'd8588344, 24'd8262247, 24'd7961156, 24'd7744657, 24'd7655595, 24'd7711594, 24'd7901574, 24'd8187936, 24'd8514011, 24'd8815269, 24'd9032091, 
24'd9121569, 24'd9065996, 24'd8876368, 24'd8590214, 24'd8264162, 24'd7962737, 24'd7745592, 24'd7655698, 24'd7710846, 24'd7900121, 24'd8186067, 24'd8512096, 24'd8813686, 24'd9031154, 24'd9121463, 24'd9066742, 24'd8877819, 24'd8592082, 24'd8266077, 24'd7964322, 24'd7746531, 24'd7655807, 24'd7710102, 24'd7898672, 24'd8184200, 24'd8510179, 24'd8812100, 24'd9030212, 24'd9121352, 24'd9067483, 
24'd8879266, 24'd8593948, 24'd8267994, 24'd7965909, 24'd7747475, 24'd7655921, 24'd7709363, 24'd7897227, 24'd8182334, 24'd8508262, 24'd8810511, 24'd9029266, 24'd9121236, 24'd9068220, 24'd8880710, 24'd8595814, 24'd8269912, 24'd7967500, 24'd7748424, 24'd7656039, 24'd7708629, 24'd7895785, 24'd8180469, 24'd8506344, 24'd8808919, 24'd9028315, 24'd9121114, 24'd9068952, 24'd8882150, 24'd8597677, 
24'd8271830, 24'd7969093, 24'd7749377, 24'd7656163, 24'd7707899, 24'd7894346, 24'd8178606, 24'd8504425, 24'd8807324, 24'd9027360, 24'd9120988, 24'd9069679, 24'd8883587, 24'd8599540, 24'd8273749, 24'd7970689, 24'd7750334, 24'd7656293, 24'd7707175, 24'd7892911, 24'd8176745, 24'd8502506, 24'd8805726, 24'd9026400, 24'd9120856, 24'd9070401, 24'd8885020, 24'd8601401, 24'd8275669, 24'd7972289, 
24'd7751296, 24'd7656427, 24'd7706455, 24'd7891479, 24'd8174885, 24'd8500585, 24'd8804126, 24'd9025436, 24'd9120719, 24'd9071118, 24'd8886450, 24'd8603260, 24'd8277590, 24'd7973891, 24'd7752263, 24'd7656566, 24'd7705740, 24'd7890051, 24'd8173026, 24'd8498664, 24'd8802522, 24'd9024467, 24'd9120577, 24'd9071831, 24'd8887877, 24'd8605118, 24'd8279512, 24'd7975496, 24'd7753234, 24'd7656711, 
24'd7705029, 24'd7888626, 24'd8171169, 24'd8496742, 24'd8800916, 24'd9023494, 24'd9120430, 24'd9072539, 24'd8889300, 24'd8606974, 24'd8281434, 24'd7977104, 24'd7754209, 24'd7656861, 24'd7704324, 24'd7887205, 24'd8169313, 24'd8494819, 24'd8799306, 24'd9022517, 24'd9120277, 24'd9073242, 24'd8890719, 24'd8608829, 24'd8283357, 24'd7978715, 24'd7755189, 24'd7657016, 24'd7703623, 24'd7885788, 
24'd8167459, 24'd8492896, 24'd8797694, 24'd9021535, 24'd9120120, 24'd9073941, 24'd8892135, 24'd8610682, 24'd8285281, 24'd7980328, 24'd7756173, 24'd7657176, 24'd7702927, 24'd7884373, 24'd8165607, 24'd8490972, 24'd8796079, 24'd9020548, 24'd9119958, 24'd9074634, 24'd8893547, 24'd8612534, 24'd8287206, 24'd7981945, 24'd7757162, 24'd7657341, 24'd7702236, 24'd7882963, 24'd8163756, 24'd8489047, 
24'd8794461, 24'd9019557, 24'd9119790, 24'd9075323, 24'd8894956, 24'd8614384, 24'd8289131, 24'd7983564, 24'd7758155, 24'd7657511, 24'd7701550, 24'd7881556, 24'd8161906, 24'd8487121, 24'd8792840, 24'd9018562, 24'd9119617, 24'd9076007, 24'd8896361, 24'd8616233, 24'd8291057, 24'd7985187, 24'd7759152, 24'd7657686, 24'd7700868, 24'd7880152, 24'd8160059, 24'd8485195, 24'd8791216, 24'd9017562, 
24'd9119439, 24'd9076686, 24'd8897763, 24'd8618080, 24'd8292984, 24'd7986812, 24'd7760154, 24'd7657867, 24'd7700191, 24'd7878752, 24'd8158213, 24'd8483268, 24'd8789590, 24'd9016558, 24'd9119256, 24'd9077360, 24'd8899161, 24'd8619925, 24'd8294911, 24'd7988440, 24'd7761161, 24'd7658052, 24'd7699519, 24'd7877356, 24'd8156368, 24'd8481340, 24'd8787960, 24'd9015549, 24'd9119068, 24'd9078030, 
24'd8900556, 24'd8621769, 24'd8296839, 24'd7990070, 24'd7762171, 24'd7658243, 24'd7698852, 24'd7875963, 24'd8154525, 24'd8479412, 24'd8786328, 24'd9014537, 24'd9118875, 24'd9078694, 24'd8901947, 24'd8623611, 24'd8298768, 24'd7991704, 24'd7763187, 24'd7658439, 24'd7698190, 24'd7874574, 24'd8152684, 24'd8477483, 24'd8784693, 24'd9013519, 24'd9118676, 24'd9079354, 24'd8903334, 24'd8625451, 
24'd8300697, 24'd7993340, 24'd7764206, 24'd7658640, 24'd7697533, 24'd7873188, 24'd8150844, 24'd8475553, 24'd8783056, 24'd9012497, 24'd9118473, 24'd9080009, 24'd8904718, 24'd8627290, 24'd8302627, 24'd7994979, 24'd7765230, 24'd7658846, 24'd7696880, 24'd7871806, 24'd8149006, 24'd8473623, 24'd8781415, 24'd9011471, 24'd9118264, 24'd9080659, 24'd8906098, 24'd8629127, 24'd8304557, 24'd7996621, 
24'd7766258, 24'd7659057, 24'd7696233, 24'd7870428, 24'd8147170, 24'd8471692, 24'd8779772, 24'd9010441, 24'd9118050, 24'd9081304, 24'd8907475, 24'd8630962, 24'd8306489, 24'd7998266, 24'd7767291, 24'd7659273, 24'd7695590, 24'd7869053, 24'd8145335, 24'd8469761, 24'd8778126, 24'd9009406, 24'd9117831, 24'd9081945, 24'd8908848, 24'd8632796, 24'd8308420, 24'd7999913, 24'd7768328, 24'd7659495, 
24'd7694952, 24'd7867682, 24'd8143503, 24'd8467829, 24'd8776477, 24'd9008367, 24'd9117607, 24'd9082580, 24'd8910217, 24'd8634628, 24'd8310352, 24'd8001563, 24'd7769369, 24'd7659721, 24'd7694319, 24'd7866315, 24'd8141671, 24'd8465896, 24'd8774826, 24'd9007323, 24'd9117378, 24'd9083211, 24'd8911583, 24'd8636458, 24'd8312285, 24'd8003216, 24'd7770415, 24'd7659953, 24'd7693691, 24'd7864951, 
24'd8139842, 24'd8463963, 24'd8773172, 24'd9006276, 24'd9117144, 24'd9083837, 24'd8912944, 24'd8638287, 24'd8314218, 24'd8004871, 24'd7771465, 24'd7660190, 24'd7693067, 24'd7863591, 24'd8138014, 24'd8462030, 24'd8771515, 24'd9005223, 24'd9116905, 24'd9084458, 24'd8914303, 24'd8640114, 24'd8316152, 24'd8006530, 24'd7772519, 24'd7660432, 24'd7692449, 24'd7862235, 24'd8136188, 24'd8460096, 
24'd8769855, 24'd9004167, 24'd9116660, 24'd9085074, 24'd8915657, 24'd8641939, 24'd8318087, 24'd8008190, 24'd7773578, 24'd7660679, 24'd7691835, 24'd7860882, 24'd8134364, 24'd8458161, 24'd8768193, 24'd9003106, 24'd9116411, 24'd9085685, 24'd8917008, 24'd8643762, 24'd8320021, 24'd8009854, 24'd7774641, 24'd7660931, 24'd7691227, 24'd7859533, 24'd8132542, 24'd8456226, 24'd8766528, 24'd9002041, 
24'd9116156, 24'd9086291, 24'd8918355, 24'd8645584, 24'd8321957, 24'd8011520, 24'd7775708, 24'd7661188, 24'd7690623, 24'd7858187, 24'd8130721, 24'd8454290, 24'd8764861, 24'd9000972, 24'd9115897, 24'd9086892, 24'd8919699, 24'd8647403, 24'd8323893, 24'd8013189, 24'd7776780, 24'd7661450, 24'd7690024, 24'd7856846, 24'd8128903, 24'd8452354, 24'd8763191, 24'd8999898, 24'd9115632, 24'd9087489, 
24'd8921039, 24'd8649221, 24'd8325829, 24'd8014860, 24'd7777856, 24'd7661718, 24'd7689430, 24'd7855508, 24'd8127086, 24'd8450418, 24'd8761518, 24'd8998820, 24'd9115362, 24'd9088080, 24'd8922374, 24'd8651037, 24'd8327765, 24'd8016534, 24'd7778936, 24'd7661990, 24'd7688841, 24'd7854174, 24'd8125271, 24'd8448481, 24'd8759843, 24'd8997738, 24'd9115087, 24'd9088667, 24'd8923707, 24'd8652851, 
24'd8329703, 24'd8018211, 24'd7780020, 24'd7662268, 24'd7688257, 24'd7852844, 24'd8123457, 24'd8446544, 24'd8758165, 24'd8996651, 24'd9114807, 24'd9089249, 24'd8925035, 24'd8654664, 24'd8331640, 24'd8019890, 24'd7781109, 24'd7662550, 24'd7687677, 24'd7851517, 24'd8121646, 24'd8444606, 24'd8756484, 24'd8995560, 24'd9114521, 24'd9089826, 24'd8926360, 24'd8656474, 24'd8333578, 24'd8021572, 
24'd7782202, 24'd7662838, 24'd7687103, 24'd7850194, 24'd8119836, 24'd8442668, 24'd8754801, 24'd8994465, 24'd9114231, 24'd9090398, 24'd8927681, 24'd8658283, 24'd8335516, 24'd8023257, 24'd7783299, 24'd7663131, 24'd7686533, 24'd7848875, 24'd8118029, 24'd8440729, 24'd8753115, 24'd8993366, 24'd9113936, 24'd9090965, 24'd8928998, 24'd8660089, 24'd8337455, 24'd8024943, 24'd7784400, 24'd7663429, 
24'd7685969, 24'd7847560, 24'd8116223, 24'd8438791, 24'd8751427, 24'd8992262, 24'd9113635, 24'd9091527, 24'd8930312, 24'd8661894, 24'd8339394, 24'd8026633, 24'd7785506, 24'd7663732, 24'd7685409, 24'd7846248, 24'd8114419, 24'd8436851, 24'd8749736, 24'd8991154, 24'd9113330, 24'd9092084, 24'd8931621, 24'd8663697, 24'd8341333, 24'd8028325, 24'd7786616, 24'd7664040, 24'd7684855, 24'd7844941, 
24'd8112617, 24'd8434912, 24'd8748043, 24'd8990042, 24'd9113019, 24'd9092636, 24'd8932927, 24'd8665498, 24'd8343273, 24'd8030020, 24'd7787730, 24'd7664353, 24'd7684305, 24'd7843637, 24'd8110817, 24'd8432972, 24'd8746347, 24'd8988926, 24'd9112703, 24'd9093183, 24'd8934229, 24'd8667297, 24'd8345213, 24'd8031717, 24'd7788849, 24'd7664671, 24'd7683760, 24'd7842337, 24'd8109019, 24'd8431032, 
24'd8744649, 24'd8987806, 24'd9112383, 24'd9093726, 24'd8935527, 24'd8669094, 24'd8347153, 24'd8033416, 24'd7789971, 24'd7664995, 24'd7683220, 24'd7841040, 24'd8107223, 24'd8429091, 24'd8742948, 24'd8986681, 24'd9112057, 24'd9094263, 24'd8936821, 24'd8670889, 24'd8349094, 24'd8035119, 24'd7791098, 24'd7665323, 24'd7682685, 24'd7839748, 24'd8105429, 24'd8427151, 24'd8741245, 24'd8985552, 
24'd9111726, 24'd9094795, 24'd8938112, 24'd8672682, 24'd8351035, 24'd8036823, 24'd7792229, 24'd7665657, 24'd7682155, 24'd7838459, 24'd8103637, 24'd8425210, 24'd8739539, 24'd8984419, 24'd9111390, 24'd9095323, 24'd8939398, 24'd8674473, 24'd8352976, 24'd8038530, 24'd7793364, 24'd7665995, 24'd7681630, 24'd7837175, 24'd8101847, 24'd8423268, 24'd8737830, 24'd8983282, 24'd9111049, 24'd9095845, 
24'd8940681, 24'd8676263, 24'd8354918, 24'd8040240, 24'd7794503, 24'd7666339, 24'd7681110, 24'd7835894, 24'd8100059, 24'd8421327, 24'd8736120, 24'd8982141, 24'd9110702, 24'd9096363, 24'd8941960, 24'd8678050, 24'd8356859, 24'd8041952, 24'd7795647, 24'd7666687, 24'd7680595, 24'd7834617, 24'd8098273, 24'd8419385, 24'd8734407, 24'd8980995, 24'd9110351, 24'd9096876, 24'd8943235, 24'd8679835, 
24'd8358801, 24'd8043666, 24'd7796794, 24'd7667041, 24'd7680085, 24'd7833344, 24'd8096489, 24'd8417443, 24'd8732691, 24'd8979845, 24'd9109995, 24'd9097383, 24'd8944506, 24'd8681618, 24'd8360743, 24'd8045383, 24'd7797946, 24'd7667400, 24'd7679580, 24'd7832075, 24'd8094707, 24'd8415501, 24'd8730973, 24'd8978692, 24'd9109634, 24'd9097886, 24'd8945773, 24'd8683399, 24'd8362685, 24'd8047102, 
24'd7799102, 24'd7667764, 24'd7679079, 24'd7830809, 24'd8092927, 24'd8413558, 24'd8729253, 24'd8977534, 24'd9109267, 24'd9098384, 24'd8947037, 24'd8685178, 24'd8364628, 24'd8048824, 24'd7800262, 24'd7668133, 24'd7678584, 24'd7829548, 24'd8091149, 24'd8411616, 24'd8727530, 24'd8976372, 24'd9108896, 24'd9098876, 24'd8948296, 24'd8686954, 24'd8366570, 24'd8050548, 24'd7801426, 24'd7668507, 
24'd7678094, 24'd7828291, 24'd8089373, 24'd8409673, 24'd8725805, 24'd8975205, 24'd9108519, 24'd9099364, 24'd8949552, 24'd8688729, 24'd8368513, 24'd8052274, 24'd7802594, 24'd7668886, 24'd7677609, 24'd7827037, 24'd8087599, 24'd8407730, 24'd8724077, 24'd8974035, 24'd9108138, 24'd9099847, 24'd8950803, 24'd8690502, 24'd8370456, 24'd8054003, 24'd7803767, 24'd7669270, 24'd7677128, 24'd7825788, 
24'd8085828, 24'd8405787, 24'd8722347, 24'd8972861, 24'd9107751, 24'd9100325, 24'd8952051, 24'd8692272, 24'd8372399, 24'd8055734, 24'd7804943, 24'd7669659, 24'd7676653, 24'd7824542, 24'd8084058, 24'd8403844, 24'd8720615, 24'd8971682, 24'd9107360, 24'd9100798, 24'd8953294, 24'd8694041, 24'd8374342, 24'd8057467, 24'd7806124, 24'd7670053, 24'd7676183, 24'd7823300, 24'd8082291, 24'd8401901, 
24'd8718880, 24'd8970499, 24'd9106963, 24'd9101265, 24'd8954534, 24'd8695807, 24'd8376286, 24'd8059203, 24'd7807308, 24'd7670452, 24'd7675718, 24'd7822063, 24'd8080526, 24'd8399958, 24'd8717144, 24'd8969313, 24'd9106561, 24'd9101728, 24'd8955770, 24'd8697571, 24'd8378229, 24'd8060941, 24'd7808497, 24'd7670856, 24'd7675257, 24'd7820829, 24'd8078763, 24'd8398014, 24'd8715404, 24'd8968122, 
24'd9106155, 24'd9102186, 24'd8957002, 24'd8699333, 24'd8380172, 24'd8062681, 24'd7809690, 24'd7671266, 24'd7674802, 24'd7819599, 24'd8077002, 24'd8396071, 24'd8713663, 24'd8966927, 24'd9105743, 24'd9102639, 24'd8958229, 24'd8701093, 24'd8382116, 24'd8064424, 24'd7810887, 24'd7671680, 24'd7674352, 24'd7818373, 24'd8075243, 24'd8394127, 24'd8711919, 24'd8965728, 24'd9105326, 24'd9103087, 
24'd8959453, 24'd8702850, 24'd8384059, 24'd8066169, 24'd7812088, 24'd7672099, 24'd7673906, 24'd7817152, 24'd8073487, 24'd8392184, 24'd8710173, 24'd8964525, 24'd9104904, 24'd9103529, 24'd8960673, 24'd8704606, 24'd8386003, 24'd8067916, 24'd7813293, 24'd7672524, 24'd7673466, 24'd7815934, 24'd8071733, 24'd8390240, 24'd8708425, 24'd8963318, 24'd9104477, 24'd9103967, 24'd8961889, 24'd8706359, 
24'd8387946, 24'd8069665, 24'd7814502, 24'd7672953, 24'd7673031, 24'd7814720, 24'd8069981, 24'd8388297, 24'd8706674, 24'd8962107, 24'd9104046, 24'd9104400, 24'd8963100, 24'd8708110, 24'd8389890, 24'd8071417, 24'd7815715, 24'd7673387, 24'd7672601, 24'd7813510, 24'd8068231, 24'd8386353, 24'd8704922, 24'd8960892, 24'd9103609, 24'd9104828, 24'd8964308, 24'd8709858, 24'd8391834, 24'd8073171, 
24'd7816932, 24'd7673827, 24'd7672175, 24'd7812305, 24'd8066483, 24'd8384410, 24'd8703167, 24'd8959673, 24'd9103167, 24'd9105250, 24'd8965512, 24'd8711605, 24'd8393777, 24'd8074927, 24'd7818153, 24'd7674271, 24'd7671755, 24'd7811103, 24'd8064738, 24'd8382466, 24'd8701410, 24'd8958450, 24'd9102720, 24'd9105668, 24'd8966711, 24'd8713349, 24'd8395721, 24'd8076685, 24'd7819378, 24'd7674720, 
24'd7671340, 24'd7809905, 24'd8062995, 24'd8380523, 24'd8699650, 24'd8957223, 24'd9102268, 24'd9106081, 24'd8967907, 24'd8715091, 24'd8397664, 24'd8078445, 24'd7820607, 24'd7675175, 24'd7670930, 24'd7808712, 24'd8061254, 24'd8378579, 24'd8697889, 24'd8955992, 24'd9101811, 24'd9106488, 24'd8969098, 24'd8716830, 24'd8399608, 24'd8080208, 24'd7821840, 24'd7675634, 24'd7670525, 24'd7807522, 
24'd8059516, 24'd8376636, 24'd8696125, 24'd8954757, 24'd9101349, 24'd9106891, 24'd8970286, 24'd8718568, 24'd8401551, 24'd8081973, 24'd7823077, 24'd7676099, 24'd7670125, 24'd7806337, 24'd8057780, 24'd8374693, 24'd8694359, 24'd8953518, 24'd9100882, 24'd9107289, 24'd8971469, 24'd8720303, 24'd8403494, 24'd8083740, 24'd7824318, 24'd7676568, 24'd7669730, 24'd7805156, 24'd8056046, 24'd8372749, 
24'd8692591, 24'd8952275, 24'd9100410, 24'd9107681, 24'd8972648, 24'd8722035, 24'd8405437, 24'd8085509, 24'd7825563, 24'd7677042, 24'd7669340, 24'd7803978, 24'd8054314, 24'd8370806, 24'd8690821, 24'd8951028, 24'd9099933, 24'd9108069, 24'd8973824, 24'd8723766, 24'd8407380, 24'd8087280, 24'd7826812, 24'd7677522, 24'd7668955, 24'd7802805, 24'd8052585, 24'd8368863, 24'd8689049, 24'd8949777, 
24'd9099452, 24'd9108451, 24'd8974995, 24'd8725493, 24'd8409323, 24'd8089053, 24'd7828064, 24'd7678006, 24'd7668575, 24'd7801636, 24'd8050858, 24'd8366921, 24'd8687274, 24'd8948523, 24'd9098965, 24'd9108828, 24'd8976162, 24'd8727219, 24'd8411266, 24'd8090829, 24'd7829321, 24'd7678496, 24'd7668200, 24'd7800471, 24'd8049134, 24'd8364978, 24'd8685498, 24'd8947264, 24'd9098473, 24'd9109201, 
24'd8977325, 24'd8728942, 24'd8413208, 24'd8092606, 24'd7830582, 24'd7678990, 24'd7667830, 24'd7799311, 24'd8047412, 24'd8363035, 24'd8683719, 24'd8946001, 24'd9097976, 24'd9109568, 24'd8978483, 24'd8730663, 24'd8415151, 24'd8094386, 24'd7831846, 24'd7679489, 24'd7667465, 24'd7798154, 24'd8045692, 24'd8361093, 24'd8681939, 24'd8944735, 24'd9097474, 24'd9109930, 24'd8979638, 24'd8732382, 
24'd8417093, 24'd8096167, 24'd7833115, 24'd7679993, 24'd7667105, 24'd7797001, 24'd8043975, 24'd8359151, 24'd8680156, 24'd8943464, 24'd9096968, 24'd9110287, 24'd8980788, 24'd8734098, 24'd8419035, 24'd8097951, 24'd7834387, 24'd7680503, 24'd7666751, 24'd7795853, 24'd8042260, 24'd8357209, 24'd8678371, 24'd8942190, 24'd9096456, 24'd9110640, 24'd8981935, 24'd8735811, 24'd8420977, 24'd8099737, 
24'd7835663, 24'd7681017, 24'd7666401, 24'd7794709, 24'd8040548, 24'd8355267, 24'd8676585, 24'd8940912, 24'd9095939, 24'd9110987, 24'd8983077, 24'd8737522, 24'd8422918, 24'd8101524, 24'd7836944, 24'd7681536, 24'd7666057, 24'd7793569, 24'd8038838, 24'd8353326, 24'd8674796, 24'd8939630, 24'd9095417, 24'd9111329, 24'd8984215, 24'd8739231, 24'd8424860, 24'd8103314, 24'd7838228, 24'd7682060, 
24'd7665717, 24'd7792433, 24'd8037131, 24'd8351385, 24'd8673005, 24'd8938344, 24'd9094891, 24'd9111666, 24'd8985348, 24'd8740937, 24'd8426801, 24'd8105106, 24'd7839515, 24'd7682589, 24'd7665383, 24'd7791301, 24'd8035425, 24'd8349444, 24'd8671212, 24'd8937054, 24'd9094359, 24'd9111997, 24'd8986478, 24'd8742641, 24'd8428742, 24'd8106900, 24'd7840807, 24'd7683123, 24'd7665054, 24'd7790174, 
24'd8033723, 24'd8347503, 24'd8669418, 24'd8935761, 24'd9093823, 24'd9112324, 24'd8987603, 24'd8744342, 24'd8430682, 24'd8108695, 24'd7842103, 24'd7683662, 24'd7664729, 24'd7789050, 24'd8032023, 24'd8345563, 24'd8667621, 24'd8934463, 24'd9093281, 24'd9112646, 24'd8988725, 24'd8746041, 24'd8432622, 24'd8110493, 24'd7843402, 24'd7684206, 24'd7664410, 24'd7787931, 24'd8030325, 24'd8343623, 
24'd8665822, 24'd8933162, 24'd9092735, 24'd9112963, 24'd8989842, 24'd8747738, 24'd8434562, 24'd8112293, 24'd7844705, 24'd7684755, 24'd7664096, 24'd7786816, 24'd8028630, 24'd8341683, 24'd8664022, 24'd8931857, 24'd9092184, 24'd9113274, 24'd8990954, 24'd8749431, 24'd8436502, 24'd8114094, 24'd7846012, 24'd7685309, 24'd7663787, 24'd7785706, 24'd8026938, 24'd8339743, 24'd8662219, 24'd8930548, 
24'd9091627, 24'd9113581, 24'd8992063, 24'd8751123, 24'd8438441, 24'd8115898, 24'd7847323, 24'd7685868, 24'd7663483, 24'd7784599, 24'd8025248, 24'd8337804, 24'd8660415, 24'd8929235, 24'd9091066, 24'd9113882, 24'd8993167, 24'd8752811, 24'd8440380, 24'd8117703, 24'd7848638, 24'd7686431, 24'd7663184, 24'd7783497, 24'd8023560, 24'd8335866, 24'd8658608, 24'd8927919, 24'd9090500, 24'd9114178, 
24'd8994267, 24'd8754497, 24'd8442319, 24'd8119510, 24'd7849956, 24'd7687000, 24'd7662891, 24'd7782399, 24'd8021875, 24'd8333927, 24'd8656800, 24'd8926598, 24'd9089929, 24'd9114469, 24'd8995363, 24'd8756181, 24'd8444257, 24'd8121320, 24'd7851278, 24'd7687573, 24'd7662602, 24'd7781305, 24'd8020193, 24'd8331989, 24'd8654990, 24'd8925274, 24'd9089353, 24'd9114756, 24'd8996455, 24'd8757862, 
24'd8446195, 24'd8123131, 24'd7852604, 24'd7688152, 24'd7662318, 24'd7780216, 24'd8018513, 24'd8330052, 24'd8653178, 24'd8923946, 24'd9088772, 24'd9115037, 24'd8997542, 24'd8759541, 24'd8448132, 24'd8124944, 24'd7853934, 24'd7688735, 24'd7662040, 24'd7779131, 24'd8016836, 24'd8328115, 24'd8651364, 24'd8922615, 24'd9088186, 24'd9115313, 24'd8998625, 24'd8761216, 24'd8450069, 24'd8126758, 
24'd7855267, 24'd7689323, 24'd7661766, 24'd7778050, 24'd8015162, 24'd8326178, 24'd8649549, 24'd8921280, 24'd9087596, 24'd9115583, 24'd8999704, 24'd8762890, 24'd8452005, 24'd8128575, 24'd7856605, 24'd7689916, 24'd7661498, 24'd7776973, 24'd8013490, 24'd8324241, 24'd8647731, 24'd8919940, 24'd9087000, 24'd9115849, 24'd9000778, 24'd8764560, 24'd8453942, 24'd8130393, 24'd7857945, 24'd7690514, 
24'd7661235, 24'd7775901, 24'd8011821, 24'd8322306, 24'd8645912, 24'd8918598, 24'd9086400, 24'd9116110, 24'd9001849, 24'd8766228, 24'd8455877, 24'd8132214, 24'd7859290, 24'd7691117, 24'd7660977, 24'd7774833, 24'd8010154, 24'd8320370, 24'd8644090, 24'd8917251, 24'd9085794, 24'd9116365, 24'd9002915, 24'd8767893, 24'd8457812, 24'd8134036, 24'd7860638, 24'd7691725, 24'd7660724, 24'd7773769, 
24'd8008490, 24'd8318435, 24'd8642268, 24'd8915901, 24'd9085184, 24'd9116616, 24'd9003976, 24'd8769556, 24'd8459747, 24'd8135860, 24'd7861990, 24'd7692338, 24'd7660476, 24'd7772710, 24'd8006829, 24'd8316501, 24'd8640443, 24'd8914547, 24'd9084569, 24'd9116861, 24'd9005033, 24'd8771216, 24'd8461681, 24'd8137685, 24'd7863346, 24'd7692956, 24'd7660233, 24'd7771655, 24'd8005170, 24'd8314567, 
24'd8638616, 24'd8913190, 24'd9083949, 24'd9117101, 24'd9006086, 24'd8772873, 24'd8463615, 24'd8139513, 24'd7864706, 24'd7693578, 24'd7659995, 24'd7770604, 24'd8003514, 24'd8312634, 24'd8636788, 24'd8911828, 24'd9083324, 24'd9117337, 24'd9007135, 24'd8774528, 24'd8465548, 24'd8141342, 24'd7866069, 24'd7694205, 24'd7659763, 24'd7769557, 24'd8001861, 24'd8310701, 24'd8634958, 24'd8910463, 
24'd9082694, 24'd9117567, 24'd9008179, 24'd8776180, 24'd8467481, 24'd8143172, 24'd7867436, 24'd7694838, 24'd7659535, 24'd7768515, 24'd8000210, 24'd8308768, 24'd8633126, 24'd8909095, 24'd9082060, 24'd9117791, 24'd9009219, 24'd8777829, 24'd8469413, 24'd8145005, 24'd7868806, 24'd7695475, 24'd7659313, 24'd7767477, 24'd7998562, 24'd8306837, 24'd8631293, 24'd8907722, 24'd9081420, 24'd9118011, 
24'd9010255, 24'd8779475, 24'd8471344, 24'd8146839, 24'd7870180, 24'd7696117, 24'd7659096, 24'd7766444, 24'd7996917, 24'd8304905, 24'd8629458, 24'd8906347, 24'd9080776, 24'd9118226, 24'd9011286, 24'd8781119, 24'd8473275, 24'd8148675, 24'd7871558, 24'd7696763, 24'd7658884, 24'd7765415, 24'd7995275, 24'd8302975, 24'd8627621, 24'd8904967, 24'd9080126, 24'd9118436, 24'd9012313, 24'd8782760, 
24'd8475205, 24'd8150513, 24'd7872939, 24'd7697415, 24'd7658677, 24'd7764390, 24'd7993635, 24'd8301045, 24'd8625783, 24'd8903584, 24'd9079472, 24'd9118640, 24'd9013335, 24'd8784398, 24'd8477135, 24'd8152352, 24'd7874324, 24'd7698071, 24'd7658475, 24'd7763370, 24'd7991999, 24'd8299115, 24'd8623942, 24'd8902197, 24'd9078814, 24'd9118839, 24'd9014354, 24'd8786034, 24'd8479064, 24'd8154193, 
24'd7875712, 24'd7698733, 24'd7658278, 24'd7762354, 24'd7990365, 24'd8297187, 24'd8622101, 24'd8900807, 24'd9078150, 24'd9119033, 24'd9015367, 24'd8787666, 24'd8480993, 24'd8156036, 24'd7877105, 24'd7699399, 24'd7658086, 24'd7761343, 24'd7988733, 24'd8295258, 24'd8620257, 24'd8899413, 24'd9077481, 24'd9119223, 24'd9016377, 24'd8789296, 24'd8482920, 24'd8157880, 24'd7878500, 24'd7700070, 
24'd7657900, 24'd7760335, 24'd7987105, 24'd8293331, 24'd8618412, 24'd8898015, 24'd9076808, 24'd9119407, 24'd9017382, 24'd8790923, 24'd8484847, 24'd8159726, 24'd7879900, 24'd7700746, 24'd7657718, 24'd7759333, 24'd7985479, 24'd8291404, 24'd8616566, 24'd8896614, 24'd9076130, 24'd9119585, 24'd9018382, 24'd8792547, 24'd8486774, 24'd8161573, 24'd7881303, 24'd7701426, 24'd7657542, 24'd7758334, 
24'd7983856, 24'd8289478, 24'd8614717, 24'd8895210, 24'd9075446, 24'd9119759, 24'd9019378, 24'd8794169, 24'd8488700, 24'd8163422, 24'd7882709, 24'd7702112, 24'd7657371, 24'd7757340, 24'd7982237, 24'd8287553, 24'd8612867, 24'd8893801, 24'd9074759, 24'd9119928, 24'd9020370, 24'd8795787, 24'd8490625, 24'd8165273, 24'd7884119, 24'd7702802, 24'd7657205, 24'd7756351, 24'd7980619, 24'd8285628, 
24'd8611016, 24'd8892390, 24'd9074066, 24'd9120091, 24'd9021357, 24'd8797403, 24'd8492549, 24'd8167125, 24'd7885532, 24'd7703497, 24'd7657044, 24'd7755366, 24'd7979005, 24'd8283704, 24'd8609163, 24'd8890974, 24'd9073368, 24'd9120250, 24'd9022340, 24'd8799016, 24'd8494473, 24'd8168979, 24'd7886949, 24'd7704197, 24'd7656888, 24'd7754385, 24'd7977394, 24'd8281781, 24'd8607308, 24'd8889556, 
24'd9072666, 24'd9120403, 24'd9023318, 24'd8800626, 24'd8496396, 24'd8170834, 24'd7888370, 24'd7704902, 24'd7656738, 24'd7753409, 24'd7975785, 24'd8279858, 24'd8605452, 24'd8888133, 24'd9071959, 24'd9120551, 24'd9024292, 24'd8802233, 24'd8498318, 24'd8172691, 24'd7889794, 24'd7705611, 24'd7656592, 24'd7752437, 24'd7974180, 24'd8277936, 24'd8603595, 24'd8886708, 24'd9071247, 24'd9120694, 
24'd9025262, 24'd8803837, 24'd8500239, 24'd8174550, 24'd7891222, 24'd7706326, 24'd7656452, 24'd7751470, 24'd7972577, 24'd8276016, 24'd8601736, 24'd8885278, 24'd9070531, 24'd9120832, 24'd9026227, 24'd8805438, 24'd8502160, 24'd8176409, 24'd7892653, 24'd7707045, 24'd7656316, 24'd7750507, 24'd7970977, 24'd8274095, 24'd8599875, 24'd8883845, 24'd9069809, 24'd9120964, 24'd9027187, 24'd8807037, 
24'd8504079, 24'd8178271, 24'd7894087, 24'd7707768, 24'd7656186, 24'd7749549, 24'd7969380, 24'd8272176, 24'd8598013, 24'd8882409, 24'd9069083, 24'd9121092, 24'd9028143, 24'd8808632, 24'd8505998, 24'd8180134, 24'd7895525, 24'd7708497, 24'd7656061, 24'd7748595, 24'd7967787, 24'd8270257, 24'd8596150, 24'd8880969, 24'd9068352, 24'd9121214, 24'd9029095, 24'd8810224, 24'd8507917, 24'd8181998, 
24'd7896967, 24'd7709230, 24'd7655942, 24'd7747646, 24'd7966196, 24'd8268340, 24'd8594285, 24'd8879526, 24'd9067616, 24'd9121331, 24'd9030042, 24'd8811814, 24'd8509834, 24'd8183863, 24'd7898412, 24'd7709969, 24'd7655827, 24'd7746701, 24'd7964608, 24'd8266423, 24'd8592418, 24'd8878080, 24'd9066876, 24'd9121444, 24'd9030985, 24'd8813400, 24'd8511750, 24'd8185731, 24'd7899860, 24'd7710711, 
24'd7655717, 24'd7745761, 24'd7963023, 24'd8264507, 24'd8590550, 24'd8876630, 24'd9066130, 24'd9121551, 24'd9031923, 24'd8814984, 24'd8513666, 24'd8187599, 24'd7901312, 24'd7711459, 24'd7655613, 24'd7744825, 24'd7961441, 24'd8262592, 24'd8588681, 24'd8875176, 24'd9065380, 24'd9121652, 24'd9032856, 24'd8816564, 24'd8515581, 24'd8189469, 24'd7902767, 24'd7712211, 24'd7655514, 24'd7743894, 
24'd7959861, 24'd8260677, 24'd8586810, 24'd8873719, 24'd9064626, 24'd9121749, 24'd9033785, 24'd8818142, 24'd8517494, 24'd8191341, 24'd7904225, 24'd7712969, 24'd7655419, 24'd7742967, 24'd7958285, 24'd8258764, 24'd8584938, 24'd8872259, 24'd9063866, 24'd9121841, 24'd9034710, 24'd8819716, 24'd8519407, 24'd8193213, 24'd7905687, 24'd7713730, 24'd7655330, 24'd7742045, 24'd7956712, 24'd8256851, 
24'd8583065, 24'd8870795, 24'd9063102, 24'd9121927, 24'd9035630, 24'd8821288, 24'd8521319, 24'd8195087, 24'd7907153, 24'd7714497, 24'd7655247, 24'd7741127, 24'd7955142, 24'd8254940, 24'd8581190, 24'd8869328, 24'd9062333, 24'd9122008, 24'd9036545, 24'd8822856, 24'd8523231, 24'd8196963, 24'd7908621, 24'd7715268, 24'd7655168, 24'd7740214, 24'd7953575, 24'd8253029, 24'd8579314, 24'd8867858, 
24'd9061559, 24'd9122085, 24'd9037456, 24'd8824422, 24'd8525141, 24'd8198840, 24'd7910094, 24'd7716044, 24'd7655094, 24'd7739305, 24'd7952012, 24'd8251120, 24'd8577436, 24'd8866384, 24'd9060781, 24'd9122156, 24'd9038363, 24'd8825984, 24'd8527050, 24'd8200718, 24'd7911569, 24'd7716825, 24'd7655026, 24'd7738401, 24'd7950451, 24'd8249211, 24'd8575557, 24'd8864907, 24'd9059998, 24'd9122221, 
24'd9039264, 24'd8827544, 24'd8528958, 24'd8202597, 24'd7913048, 24'd7717611, 24'd7654963, 24'd7737501, 24'd7948893, 24'd8247303, 24'd8573677, 24'd8863426, 24'd9059210, 24'd9122282, 24'd9040162, 24'd8829100, 24'd8530865, 24'd8204478, 24'd7914530, 24'd7718401, 24'd7654904, 24'd7736606, 24'd7947338, 24'd8245397, 24'd8571796, 24'd8861943, 24'd9058417, 24'd9122338, 24'd9041054, 24'd8830653, 
24'd8532771, 24'd8206360, 24'd7916015, 24'd7719196, 24'd7654851, 24'd7735716, 24'd7945787, 24'd8243491, 24'd8569913, 24'd8860456, 24'd9057620, 24'd9122388, 24'd9041942, 24'd8832203, 24'd8534677, 24'd8208244, 24'd7917504, 24'd7719995, 24'd7654804, 24'd7734830, 24'd7944238, 24'd8241586, 24'd8568029, 24'd8858965, 24'd9056818, 24'd9122433, 24'd9042826, 24'd8833750, 24'd8536581, 24'd8210128, 
24'd7918996, 24'd7720800, 24'd7654761, 24'd7733949, 24'd7942693, 24'd8239682, 24'd8566144, 24'd8857471, 24'd9056011, 24'd9122474, 24'd9043705, 24'd8835294, 24'd8538484, 24'd8212014, 24'd7920492, 24'd7721609, 24'd7654723, 24'd7733072, 24'd7941151, 24'd8237780, 24'd8564257, 24'd8855974, 24'd9055200, 24'd9122509, 24'd9044579, 24'd8836834, 24'd8540386, 24'd8213901, 24'd7921990, 24'd7722422, 
24'd7654691, 24'd7732200, 24'd7939612, 24'd8235878, 24'd8562370, 24'd8854474, 24'd9054384, 24'd9122538, 24'd9045449, 24'd8838372, 24'd8542287, 24'd8215790, 24'd7923492, 24'd7723240, 24'd7654664, 24'd7731333, 24'd7938076, 24'd8233978, 24'd8560481, 24'd8852971, 24'd9053564, 24'd9122563, 24'd9046314, 24'd8839906, 24'd8544187, 24'd8217679, 24'd7924997, 24'd7724063, 24'd7654641, 24'd7730470, 
24'd7936543, 24'd8232078, 24'd8558591, 24'd8851464, 24'd9052738, 24'd9122583, 24'd9047175, 24'd8841437, 24'd8546086, 24'd8219570, 24'd7926506, 24'd7724891, 24'd7654624, 24'd7729612, 24'd7935013, 24'd8230180, 24'd8556699, 24'd8849954, 24'd9051908, 24'd9122597, 24'd9048031, 24'd8842965, 24'd8547984, 24'd8221462, 24'd7928018, 24'd7725723, 24'd7654613, 24'd7728758, 24'd7933487, 24'd8228283, 
24'd8554807, 24'd8848440, 24'd9051074, 24'd9122606, 24'd9048882, 24'd8844490, 24'd8549880, 24'd8223355, 24'd7929533, 24'd7726560, 24'd7654606, 24'd7727909, 24'd7931963, 24'd8226387, 24'd8552913, 24'd8846924, 24'd9050235, 24'd9122610, 24'd9049729, 24'd8846012, 24'd8551776, 24'd8225249, 24'd7931051, 24'd7727402, 24'd7654604, 24'd7727065, 24'd7930443, 24'd8224492, 24'd8551018, 24'd8845404, 
24'd9049391, 24'd9122609, 24'd9050571, 24'd8847530, 24'd8553670, 24'd8227145, 24'd7932572, 24'd7728248, 24'd7654608, 24'd7726225, 24'd7928927, 24'd8222598, 24'd8549122, 24'd8843881, 24'd9048542, 24'd9122603, 24'd9051408, 24'd8849046, 24'd8555564, 24'd8229041, 24'd7934097, 24'd7729099, 24'd7654617, 24'd7725390, 24'd7927413, 24'd8220705, 24'd8547225, 24'd8842355, 24'd9047689, 24'd9122592, 
24'd9052241, 24'd8850558, 24'd8557456, 24'd8230939, 24'd7935624, 24'd7729954, 24'd7654631, 24'd7724560, 24'd7925903, 24'd8218814, 24'd8545327, 24'd8840826, 24'd9046831, 24'd9122575, 24'd9053069, 24'd8852066, 24'd8559346, 24'd8232837, 24'd7937155, 24'd7730814, 24'd7654650, 24'd7723734, 24'd7924395, 24'd8216924, 24'd8543428, 24'd8839293, 24'd9045969, 24'd9122554, 24'd9053892, 24'd8853572, 
24'd8561236, 24'd8234737, 24'd7938689, 24'd7731679, 24'd7654674, 24'd7722913, 24'd7922892, 24'd8215035, 24'd8541527, 24'd8837758, 24'd9045102, 24'd9122527, 24'd9054711, 24'd8855074, 24'd8563125, 24'd8236638, 24'd7940226, 24'd7732548, 24'd7654703, 24'd7722096, 24'd7921391, 24'd8213147, 24'd8539626, 24'd8836219, 24'd9044230, 24'd9122495, 24'd9055525, 24'd8856573, 24'd8565012, 24'd8238540, 
24'd7941767, 24'd7733422, 24'd7654738, 24'd7721285, 24'd7919894, 24'd8211260, 24'd8537723, 24'd8834677, 24'd9043354, 24'd9122458, 24'd9056334, 24'd8858069, 24'd8566898, 24'd8240443, 24'd7943310, 24'd7734301, 24'd7654777, 24'd7720478, 24'd7918399, 24'd8209375, 24'd8535820, 24'd8833132, 24'd9042473, 24'd9122416, 24'd9057139, 24'd8859561, 24'd8568782, 24'd8242347, 24'd7944857, 24'd7735184, 
24'd7654822, 24'd7719675, 24'd7916909, 24'd8207491, 24'd8533915, 24'd8831584, 24'd9041588, 24'd9122369, 24'd9057939, 24'd8861050, 24'd8570666, 24'd8244252, 24'd7946407, 24'd7736071, 24'd7654872, 24'd7718877, 24'd7915421, 24'd8205608, 24'd8532010, 24'd8830032, 24'd9040698, 24'd9122316, 24'd9058735, 24'd8862536, 24'd8572548, 24'd8246159, 24'd7947959, 24'd7736964, 24'd7654927, 24'd7718084, 
24'd7913937, 24'd8203726, 24'd8530103, 24'd8828478, 24'd9039803, 24'd9122258, 24'd9059525, 24'd8864019, 24'd8574429, 24'd8248066, 24'd7949515, 24'd7737860, 24'd7654987, 24'd7717296, 24'd7912456, 24'd8201846, 24'd8528195, 24'd8826921, 24'd9038904, 24'd9122196, 24'd9060311, 24'd8865498, 24'd8576309, 24'd8249974, 24'd7951074, 24'd7738762, 24'd7655053, 24'd7716513, 24'd7910979, 24'd8199967, 
24'd8526287, 24'd8825360, 24'd9038001, 24'd9122128, 24'd9061092, 24'd8866974, 24'd8578187, 24'd8251883, 24'd7952636, 24'd7739668, 24'd7655123, 24'd7715734, 24'd7909505, 24'd8198089, 24'd8524377, 24'd8823796, 24'd9037093, 24'd9122055, 24'd9061869, 24'd8868446, 24'd8580064, 24'd8253793, 24'd7954202, 24'd7740578, 24'd7655199, 24'd7714959, 24'd7908034, 24'd8196213, 24'd8522467, 24'd8822230, 
24'd9036180, 24'd9121977, 24'd9062641, 24'd8869915, 24'd8581940, 24'd8255704, 24'd7955770, 24'd7741493, 24'd7655280, 24'd7714190, 24'd7906567, 24'd8194338, 24'd8520555, 24'd8820660, 24'd9035263, 24'd9121893, 24'd9063408, 24'd8871381, 24'd8583814, 24'd8257616, 24'd7957341, 24'd7742413, 24'd7655365, 24'd7713425, 24'd7905103, 24'd8192465, 24'd8518643, 24'd8819087, 24'd9034341, 24'd9121805, 
24'd9064170, 24'd8872843, 24'd8585687, 24'd8259529, 24'd7958915, 24'd7743337, 24'd7655456, 24'd7712665, 24'd7903642, 24'd8190592, 24'd8516730, 24'd8817512, 24'd9033414, 24'd9121711, 24'd9064928, 24'd8874302, 24'd8587558, 24'd8261442, 24'd7960492, 24'd7744265, 24'd7655553, 24'd7711910, 24'd7902185, 24'd8188722, 24'd8514815, 24'd8815933, 24'd9032484, 24'd9121612, 24'd9065681, 24'd8875758, 
24'd8589428, 24'd8263357, 24'd7962073, 24'd7745199, 24'd7655654, 24'd7711160, 24'd7900731, 24'd8186852, 24'd8512900, 24'd8814351, 24'd9031548, 24'd9121508, 24'd9066429, 24'd8877210, 24'd8591297, 24'd8265273, 24'd7963656, 24'd7746136, 24'd7655760, 24'd7710414, 24'd7899281, 24'd8184984, 24'd8510984, 24'd8812766, 24'd9030608, 24'd9121399, 24'd9067172, 24'd8878658, 24'd8593164, 24'd8267189, 
24'd7965242, 24'd7747078, 24'd7655872, 24'd7709673, 24'd7897834, 24'd8183118, 24'd8509068, 24'd8811179, 24'd9029664, 24'd9121285, 24'd9067911, 24'd8880104, 24'd8595030, 24'd8269106, 24'd7966831, 24'd7748025, 24'd7655989, 24'd7708937, 24'd7896390, 24'd8181252, 24'd8507150, 24'd8809588, 24'd9028715, 24'd9121166, 24'd9068645, 24'd8881545, 24'd8596895, 24'd8271024, 24'd7968423, 24'd7748976, 
24'd7656111, 24'd7708205, 24'd7894950, 24'd8179389, 24'd8505231, 24'd8807995, 24'd9027762, 24'd9121041, 24'd9069374, 24'd8882984, 24'd8598758, 24'd8272943, 24'd7970018, 24'd7749932, 24'd7656238, 24'd7707478, 24'd7893513, 24'd8177526, 24'd8503312, 24'd8806398, 24'd9026804, 24'd9120912, 24'd9070098, 24'd8884419, 24'd8600619, 24'd8274863, 24'd7971616, 24'd7750892, 24'd7656370, 24'd7706757, 
24'd7892080, 24'd8175666, 24'd8501392, 24'd8804798, 24'd9025841, 24'd9120777, 24'd9070818, 24'd8885850, 24'd8602479, 24'd8276783, 24'd7973217, 24'd7751856, 24'd7656507, 24'd7706039, 24'd7890651, 24'd8173806, 24'd8499471, 24'd8803196, 24'd9024875, 24'd9120637, 24'd9071532, 24'd8887278, 24'd8604338, 24'd8278705, 24'd7974821, 24'd7752825, 24'd7656650, 24'd7705327, 24'd7889224, 24'd8171949, 
24'd8497549, 24'd8801591, 24'd9023903, 24'd9120492, 24'd9072242, 24'd8888702, 24'd8606195, 24'd8280627, 24'd7976428, 24'd7753799, 24'd7656797, 24'd7704619, 24'd7887802, 24'd8170093, 24'd8495627, 24'd8799983, 24'd9022928, 24'd9120342, 24'd9072947, 24'd8890123, 24'd8608050, 24'd8282549, 24'd7978038, 24'd7754777, 24'd7656950, 24'd7703917, 24'd7886383, 24'd8168238, 24'd8493704, 24'd8798371, 
24'd9021948, 24'd9120187, 24'd9073648, 24'd8891541, 24'd8609904, 24'd8284473, 24'd7979650, 24'd7755759, 24'd7657108, 24'd7703219, 24'd7884967, 24'd8166385, 24'd8491780, 24'd8796758, 24'd9020963, 24'd9120026, 24'd9074343, 24'd8892955, 24'd8611756, 24'd8286397, 24'd7981266, 24'd7756746, 24'd7657271, 24'd7702526, 24'd7883555, 24'd8164533, 24'd8489855, 24'd8795141, 24'd9019974, 24'd9119861, 
24'd9075034, 24'd8894365, 24'd8613607, 24'd8288322, 24'd7982884, 24'd7757737, 24'd7657439, 24'd7701837, 24'd7882146, 24'd8162683, 24'd8487930, 24'd8793521, 24'd9018981, 24'd9119690, 24'd9075720, 24'd8895772, 24'd8615456, 24'd8290248, 24'd7984505, 24'd7758733, 24'd7657612, 24'd7701154, 24'd7880741, 24'd8160835, 24'd8486004, 24'd8791899, 24'd9017983, 24'd9119515, 24'd9076401, 24'd8897175, 
24'd8617304, 24'd8292174, 24'd7986129, 24'd7759733, 24'd7657790, 24'd7700475, 24'd7879340, 24'd8158988, 24'd8484077, 24'd8790273, 24'd9016980, 24'd9119334, 24'd9077078, 24'd8898575, 24'd8619150, 24'd8294101, 24'd7987756, 24'd7760737, 24'd7657974, 24'd7699801, 24'd7877942, 24'd8157143, 24'd8482150, 24'd8788645, 24'd9015974, 24'd9119148, 24'd9077749, 24'd8899971, 24'd8620994, 24'd8296029, 
24'd7989385, 24'd7761746, 24'd7658162, 24'd7699132, 24'd7876548, 24'd8155299, 24'd8480222, 24'd8787014, 24'd9014963, 24'd9118956, 24'd9078416, 24'd8901363, 24'd8622837, 24'd8297958, 24'd7991017, 24'd7762760, 24'd7658356, 24'd7698468, 24'd7875157, 24'd8153457, 24'd8478293, 24'd8785380, 24'd9013947, 24'd9118760, 24'd9079077, 24'd8902752, 24'd8624678, 24'd8299887, 24'd7992653, 24'd7763777, 
24'd7658555, 24'd7697808, 24'd7873770, 24'd8151617, 24'd8476364, 24'd8783744, 24'd9012927, 24'd9118559, 24'd9079734, 24'd8904137, 24'd8626518, 24'd8301816, 24'd7994290, 24'd7764799, 24'd7658759, 24'd7697154, 24'd7872386, 24'd8149778, 24'd8474434, 24'd8782105, 24'd9011903, 24'd9118352, 24'd9080387, 24'd8905519, 24'd8628356, 24'd8303746, 24'd7995931, 24'd7765826, 24'd7658968, 24'd7696504, 
24'd7871007, 24'd8147941, 24'd8472503, 24'd8780462, 24'd9010874, 24'd9118141, 24'd9081034, 24'd8906897, 24'd8630192, 24'd8305677, 24'd7997575, 24'd7766857, 24'd7659182, 24'd7695859, 24'd7869630, 24'd8146106, 24'd8470572, 24'd8778818, 24'd9009841, 24'd9117924, 24'd9081676, 24'd8908271, 24'd8632026, 24'd8307609, 24'd7999221, 24'd7767892, 24'd7659401, 24'd7695219, 24'd7868258, 24'd8144272, 
24'd8468640, 24'd8777170, 24'd9008804, 24'd9117702, 24'd9082314, 24'd8909642, 24'd8633859, 24'd8309541, 24'd8000870, 24'd7768931, 24'd7659626, 24'd7694584, 24'd7866889, 24'd8142440, 24'd8466708, 24'd8775520, 24'd9007762, 24'd9117475, 24'd9082947, 24'd8911009, 24'd8635690, 24'd8311473, 24'd8002521, 24'd7769975, 24'd7659855, 24'd7693954, 24'd7865523, 24'd8140610, 24'd8464775, 24'd8773867, 
24'd9006716, 24'd9117243, 24'd9083574, 24'd8912373, 24'd8637519, 24'd8313406, 24'd8004176, 24'd7771023, 24'd7660090, 24'd7693329, 24'd7864162, 24'd8138782, 24'd8462842, 24'd8772211, 24'd9005666, 24'd9117006, 24'd9084197, 24'd8913733, 24'd8639347, 24'd8315340, 24'd8005833, 24'd7772076, 24'd7660330, 24'd7692708, 24'd7862804, 24'd8136955, 24'd8460908, 24'd8770553, 24'd9004611, 24'd9116764, 
24'd9084815, 24'd8915089, 24'd8641172, 24'd8317274, 24'd8007492, 24'd7773133, 24'd7660574, 24'd7692092, 24'd7861450, 24'd8135130, 24'd8458974, 24'd8768892, 24'd9003552, 24'd9116516, 24'd9085429, 24'd8916441, 24'd8642996, 24'd8319209, 24'd8009155, 24'd7774194, 24'd7660824, 24'd7691482, 24'd7860099, 24'd8133307, 24'd8457039, 24'd8767228, 24'd9002489, 24'd9116264, 24'd9086037, 24'd8917790, 
24'd8644819, 24'd8321144, 24'd8010820, 24'd7775259, 24'd7661079, 24'd7690876, 24'd7858752, 24'd8131486, 24'd8455103, 24'd8765562, 24'd9001421, 24'd9116006, 24'd9086640, 24'd8919135, 24'd8646639, 24'd8323079, 24'd8012488, 24'd7776329, 24'd7661339, 24'd7690275, 24'd7857409, 24'd8129666, 24'd8453168, 24'd8763893, 24'd9000349, 24'd9115744, 24'd9087239, 24'd8920476, 24'd8648458, 24'd8325015, 
24'd8014158, 24'd7777403, 24'd7661605, 24'd7689679, 24'd7856070, 24'd8127849, 24'd8451231, 24'd8762221, 24'd8999273, 24'd9115476, 24'd9087832, 24'd8921814, 24'd8650275, 24'd8326952, 24'd8015831, 24'd7778482, 24'd7661875, 24'd7689088, 24'd7854734, 24'd8126033, 24'd8449295, 24'd8760547, 24'd8998193, 24'd9115203, 24'd9088421, 24'd8923148, 24'd8652090, 24'd8328889, 24'd8017506, 24'd7779564, 
24'd7662150, 24'd7688501, 24'd7853402, 24'd8124219, 24'd8447358, 24'd8758870, 24'd8997108, 24'd9114925, 24'd9089005, 24'd8924478, 24'd8653903, 24'd8330826, 24'd8019185, 24'd7780651, 24'd7662431, 24'd7687920, 24'd7852074, 24'd8122407, 24'd8445420, 24'd8757190, 24'd8996019, 24'd9114642, 24'd9089584, 24'd8925804, 24'd8655714, 24'd8332764, 24'd8020865, 24'd7781742, 24'd7662717, 24'd7687344, 
24'd7850749, 24'd8120596, 24'd8443482, 24'd8755508, 24'd8994926, 24'd9114354, 24'd9090158, 24'd8927127, 24'd8657523, 24'd8334702, 24'd8022549, 24'd7782838, 24'd7663007, 24'd7686772, 24'd7849429, 24'd8118788, 24'd8441544, 24'd8753824, 24'd8993828, 24'd9114060, 24'd9090727, 24'd8928445, 24'd8659331, 24'd8336641, 24'd8024235, 24'd7783937, 24'd7663303, 24'd7686205, 24'd7848112, 24'd8116981, 
24'd8439605, 24'd8752137, 24'd8992726, 24'd9113762, 24'd9091291, 24'd8929760, 24'd8661136, 24'd8338579, 24'd8025923, 24'd7785041, 24'd7663604, 24'd7685644, 24'd7846799, 24'd8115177, 24'd8437666, 24'd8750447, 24'd8991620, 24'd9113459, 24'd9091850, 24'd8931071, 24'd8662940, 24'd8340519, 24'd8027614, 24'd7786149, 24'd7663910, 24'd7685087, 24'd7845489, 24'd8113374, 24'd8435727, 24'd8748755, 
24'd8990510, 24'd9113150, 24'd9092405, 24'd8932379, 24'd8664742, 24'd8342458, 24'd8029308, 24'd7787262, 24'd7664221, 24'd7684535, 24'd7844184, 24'd8111573, 24'd8433787, 24'd8747060, 24'd8989396, 24'd9112837, 24'd9092954, 24'd8933682, 24'd8666542, 24'd8344398, 24'd8031004, 24'd7788378, 24'd7664537, 24'd7683988, 24'd7842882, 24'd8109774, 24'd8431847, 24'd8745362, 24'd8988277, 24'd9112518, 
24'd9093498, 24'd8934982, 24'd8668340, 24'd8346338, 24'd8032702, 24'd7789499, 24'd7664858, 24'd7683446, 24'd7841584, 24'd8107977, 24'd8429906, 24'd8743663, 24'd8987154, 24'd9112194, 24'd9094038, 24'd8936278, 24'd8670135, 24'd8348279, 24'd8034403, 24'd7790624, 24'd7665185, 24'd7682909, 24'd7840290, 24'd8106182, 24'd8427966, 24'd8741960, 24'd8986027, 24'd9111865, 24'd9094572, 24'd8937570, 
24'd8671929, 24'd8350220, 24'd8036107, 24'd7791753, 24'd7665516, 24'd7682377, 24'd7839000, 24'd8104389, 24'd8426025, 24'd8740256, 24'd8984896, 24'd9111531, 24'd9095102, 24'd8938858, 24'd8673721, 24'd8352161, 24'd8037813, 24'd7792887, 24'd7665852, 24'd7681850, 24'd7837714, 24'd8102598, 24'd8424084, 24'd8738548, 24'd8983760, 24'd9111193, 24'd9095627, 24'd8940143, 24'd8675511, 24'd8354102, 
24'd8039521, 24'd7794024, 24'd7666194, 24'd7681328, 24'd7836431, 24'd8100809, 24'd8422142, 24'd8736839, 24'd8982621, 24'd9110849, 24'd9096146, 24'd8941423, 24'd8677299, 24'd8356044, 24'd8041232, 24'd7795166, 24'd7666540, 24'd7680811, 24'd7835153, 24'd8099023, 24'd8420201, 24'd8735126, 24'd8981477, 24'd9110499, 24'd9096661, 24'd8942700, 24'd8679085, 24'd8357985, 24'd8042946, 24'd7796312, 
24'd7666892, 24'd7680299, 24'd7833878, 24'd8097238, 24'd8418259, 24'd8733412, 24'd8980329, 24'd9110145, 24'd9097171, 24'd8943973, 24'd8680869, 24'd8359927, 24'd8044661, 24'd7797462, 24'd7667249, 24'd7679791, 24'd7832607, 24'd8095455, 24'd8416317, 24'd8731695, 24'd8979177, 24'd9109786, 24'd9097675, 24'd8945242, 24'd8682651, 24'd8361869, 24'd8046380, 24'd7798616, 24'd7667610, 24'd7679289, 
24'd7831340, 24'd8093674, 24'd8414374, 24'd8729975, 24'd8978021, 24'd9109422, 24'd9098175, 24'd8946507, 24'd8684431, 24'd8363812, 24'd8048100, 24'd7799774, 24'd7667977, 24'd7678792, 24'd7830077, 24'd8091895, 24'd8412432, 24'd8728254, 24'd8976860, 24'd9109053, 24'd9098670, 24'd8947768, 24'd8686208, 24'd8365754, 24'd8049823, 24'd7800937, 24'd7668349, 24'd7678299, 24'd7828818, 24'd8090119, 
24'd8410489, 24'd8726530, 24'd8975696, 24'd9108678, 24'd9099160, 24'd8949025, 24'd8687984, 24'd8367697, 24'd8051548, 24'd7802103, 24'd7668726, 24'd7677812, 24'd7827563, 24'd8088344, 24'd8408546, 24'd8724803, 24'd8974527, 24'd9108299, 24'd9099645, 24'd8950278, 24'd8689757, 24'd8369640, 24'd8053276, 24'd7803274, 24'd7669108, 24'd7677330, 24'd7826312, 24'd8086572, 24'd8406604, 24'd8723074, 
24'd8973354, 24'd9107914, 24'd9100125, 24'd8951527, 24'd8691529, 24'd8371583, 24'd8055006, 24'd7804449, 24'd7669495, 24'd7676852, 24'd7825065, 24'd8084801, 24'd8404660, 24'd8721343, 24'd8972178, 24'd9107525, 24'd9100600, 24'd8952772, 24'd8693298, 24'd8373526, 24'd8056739, 24'd7805627, 24'd7669887, 24'd7676380, 24'd7823821, 24'd8083033, 24'd8402717, 24'd8719609, 24'd8970997, 24'd9107130, 
24'd9101070, 24'd8954014, 24'd8695065, 24'd8375469, 24'd8058473, 24'd7806810, 24'd7670284, 24'd7675912, 24'd7822582, 24'd8081267, 24'd8400774, 24'd8717873, 24'd8969812, 24'd9106731, 24'd9101534, 24'd8955251, 24'd8696830, 24'd8377413, 24'd8060210, 24'd7807997, 24'd7670686, 24'd7675450, 24'd7821347, 24'd8079503, 24'd8398831, 24'd8716135, 24'd8968623, 24'd9106326, 24'd9101994, 24'd8956485, 
24'd8698593, 24'd8379356, 24'd8061950, 24'd7809188, 24'd7671093, 24'd7674993, 24'd7820115, 24'd8077741, 24'd8396887, 24'd8714395, 24'd8967429, 24'd9105916, 24'd9102449, 24'd8957714, 24'd8700354, 24'd8381299, 24'd8063691, 24'd7810384, 24'd7671505, 24'd7674540, 24'd7818888, 24'd8075982, 24'd8394944, 24'd8712652, 24'd8966232, 24'd9105502, 24'd9102899, 24'd8958940, 24'd8702112, 24'd8383243, 
24'd8065435, 24'd7811583, 24'd7671923, 24'd7674093, 24'd7817664, 24'd8074224, 24'd8393000, 24'd8710907, 24'd8965031, 24'd9105082, 24'd9103344, 24'd8960161, 24'd8703869, 24'd8385187, 24'd8067182, 24'd7812786, 24'd7672345, 24'd7673650, 24'd7816445, 24'd8072469, 24'd8391057, 24'd8709160, 24'd8963826, 24'd9104657, 24'd9103784, 24'd8961378, 24'd8705623, 24'd8387130, 24'd8068930, 24'd7813993, 
24'd7672772, 24'd7673213, 24'd7815229, 24'd8070716, 24'd8389113, 24'd8707410, 24'd8962616, 24'd9104228, 24'd9104219, 24'd8962592, 24'd8707374, 24'd8389074, 24'd8070681, 24'd7815205, 24'd7673204, 24'd7672781, 24'd7814018, 24'd8068965, 24'd8387170, 24'd8705658, 24'd8961403, 24'd9103793, 24'd9104649, 24'd8963801, 24'd8709124, 24'd8391017, 24'd8072434, 24'd7816420, 24'd7673641, 24'd7672353, 
24'd7812811, 24'd8067217, 24'd8385226, 24'd8703904, 24'd8960186, 24'd9103353, 24'd9105073, 24'd8965007, 24'd8710871, 24'd8392961, 24'd8074189, 24'd7817639, 24'd7674084, 24'd7671931, 24'd7811607, 24'd8065471, 24'd8383282, 24'd8702148, 24'd8958964, 24'd9102908, 24'd9105493, 24'd8966208, 24'd8712617, 24'd8394904, 24'd8075946, 24'd7818863, 24'd7674531, 24'd7671514, 24'd7810408, 24'd8063727, 
24'd8381339, 24'd8700390, 24'd8957739, 24'd9102458, 24'd9105908, 24'd8967405, 24'd8714359, 24'd8396848, 24'd8077706, 24'd7820090, 24'd7674983, 24'd7671101, 24'd7809213, 24'd8061985, 24'd8379395, 24'd8698629, 24'd8956510, 24'd9102004, 24'd9106318, 24'd8968598, 24'd8716100, 24'd8398791, 24'd8079467, 24'd7821322, 24'd7675441, 24'd7670694, 24'd7808022, 24'd8060246, 24'd8377452, 24'd8696866, 
24'd8955276, 24'd9101544, 24'd9106722, 24'd8969788, 24'd8717838, 24'd8400735, 24'd8081231, 24'd7822557, 24'd7675903, 24'd7670292, 24'd7806834, 24'd8058509, 24'd8375509, 24'd8695101, 24'd8954039, 24'd9101079, 24'd9107122, 24'd8970973, 24'd8719574, 24'd8402678, 24'd8082997, 24'd7823796, 24'd7676370, 24'd7669895, 24'd7805651, 24'd8056774, 24'd8373566, 24'd8693334, 24'd8952798, 24'd9100609, 
24'd9107517, 24'd8972154, 24'd8721308, 24'd8404621, 24'd8084765, 24'd7825039, 24'd7676843, 24'd7669503, 24'd7804472, 24'd8055041, 24'd8371622, 24'd8691565, 24'd8951553, 24'd9100134, 24'd9107906, 24'd8973331, 24'd8723039, 24'd8406564, 24'd8086536, 24'd7826287, 24'd7677320, 24'd7669116, 24'd7803298, 24'd8053311, 24'd8369679, 24'd8689793, 24'd8950303, 24'd9099655, 24'd9108291, 24'd8974503, 
24'd8724768, 24'd8408507, 24'd8088308, 24'd7827538, 24'd7677802, 24'd7668734, 24'd7802127, 24'd8051583, 24'd8367737, 24'd8688020, 24'd8949050, 24'd9099170, 24'd9108670, 24'd8975672, 24'd8726495, 24'd8410450, 24'd8090083, 24'd7828793, 24'd7678289, 24'd7668357, 24'd7800960, 24'd8049858, 24'd8365794, 24'd8686244, 24'd8947793, 24'd9098680, 24'd9109045, 24'd8976837, 24'd8728219, 24'd8412392, 
24'd8091859, 24'd7830052, 24'd7678782, 24'd7667985, 24'd7799798, 24'd8048135, 24'd8363851, 24'd8684467, 24'd8946532, 24'd9098185, 24'd9109414, 24'd8977997, 24'd8729941, 24'd8414335, 24'd8093638, 24'd7831315, 24'd7679279, 24'd7667618, 24'd7798639, 24'd8046414, 24'd8361909, 24'd8682687, 24'd8945267, 24'd9097686, 24'd9109779, 24'd8979153, 24'd8731660, 24'd8416277, 24'd8095419, 24'd7832582, 
24'd7679781, 24'd7667256, 24'd7797485, 24'd8044696, 24'd8359967, 24'd8680905, 24'd8943999, 24'd9097181, 24'd9110138, 24'd8980306, 24'd8733377, 24'd8418219, 24'd8097201, 24'd7833852, 24'd7680288, 24'd7666899, 24'd7796335, 24'd8042980, 24'd8358025, 24'd8679121, 24'd8942726, 24'd9096671, 24'd9110492, 24'd8981454, 24'd8735092, 24'd8420161, 24'd8098986, 24'd7835127, 24'd7680800, 24'd7666547, 
24'd7795189, 24'd8041267, 24'd8356083, 24'd8677336, 24'd8941449, 24'd9096157, 24'd9110841, 24'd8982597, 24'd8736804, 24'd8422103, 24'd8100773, 24'd7836405, 24'd7681317, 24'd7666201, 24'd7794047, 24'd8039556, 24'd8354141, 24'd8675548, 24'd8940169, 24'd9095637, 24'd9111186, 24'd8983737, 24'd8738514, 24'd8424044, 24'd8102562, 24'd7837688, 24'd7681839, 24'd7665859, 24'd7792910, 24'd8037847, 
24'd8352200, 24'd8673758, 24'd8938885, 24'd9095113, 24'd9111525, 24'd8984873, 24'd8740221, 24'd8425985, 24'd8104353, 24'd7838974, 24'd7682366, 24'd7665523, 24'd7791776, 24'd8036141, 24'd8350259, 24'd8671966, 24'd8937596, 24'd9094583, 24'd9111859, 24'd8986004, 24'd8741926, 24'd8427926, 24'd8106146, 24'd7840264, 24'd7682898, 24'd7665191, 24'd7790647, 24'd8034438, 24'd8348318, 24'd8670172, 
24'd8936304, 24'd9094049, 24'd9112188, 24'd8987131, 24'd8743628, 24'd8429867, 24'd8107941, 24'd7841558, 24'd7683435, 24'd7664865, 24'd7789522, 24'd8032737, 24'd8346378, 24'd8668376, 24'd8935009, 24'd9093509, 24'd9112511, 24'd8988254, 24'd8745328, 24'd8431807, 24'd8109738, 24'd7842856, 24'd7683977, 24'd7664544, 24'd7788401, 24'd8031038, 24'd8344438, 24'd8666578, 24'd8933709, 24'd9092965, 
24'd9112830, 24'd8989373, 24'd8747025, 24'd8433747, 24'd8111536, 24'd7844157, 24'd7684524, 24'd7664227, 24'd7787284, 24'd8029342, 24'd8342498, 24'd8664778, 24'd8932405, 24'd9092416, 24'd9113144, 24'd8990487, 24'd8748720, 24'd8435687, 24'd8113337, 24'd7845463, 24'd7685076, 24'd7663916, 24'd7786172, 24'd8027648, 24'd8340558, 24'd8662977, 24'd8931098, 24'd9091862, 24'd9113452, 24'd8991598, 
24'd8750412, 24'd8437627, 24'd8115140, 24'd7846772, 24'd7685632, 24'd7663610, 24'd7785064, 24'd8025957, 24'd8338619, 24'd8661173, 24'd8929787, 24'd9091302, 24'd9113756, 24'd8992704, 24'd8752102, 24'd8439566, 24'd8116945, 24'd7848085, 24'd7686194, 24'd7663309, 24'd7783960, 24'd8024269, 24'd8336680, 24'd8659367, 24'd8928472, 24'd9090738, 24'd9114054, 24'd8993806, 24'd8753789, 24'd8441504, 
24'd8118751, 24'd7849402, 24'd7686760, 24'd7663013, 24'd7782860, 24'd8022583, 24'd8334741, 24'd8657560, 24'd8927153, 24'd9090169, 24'd9114348, 24'd8994903, 24'd8755474, 24'd8443443, 24'd8120559, 24'd7850722, 24'd7687332, 24'd7662722, 24'd7781764, 24'd8020899, 24'd8332803, 24'd8655751, 24'd8925831, 24'd9089596, 24'd9114636, 24'd8995997, 24'd8757156, 24'd8445381, 24'd8122370, 24'd7852047, 
24'd7687908, 24'd7662437, 24'd7780673, 24'd8019219, 24'd8330866, 24'd8653939, 24'd8924505, 24'd9089017, 24'd9114919, 24'd8997086, 24'd8758836, 24'd8447318, 24'd8124182, 24'd7853375, 24'd7688489, 24'd7662156, 24'd7779586, 24'd8017540, 24'd8328928, 24'd8652126, 24'd8923175, 24'd9088433, 24'd9115197, 24'd8998171, 24'd8760513, 24'd8449255, 24'd8125996, 24'd7854707, 24'd7689076, 24'd7661881, 
24'd7778503, 24'd8015865, 24'd8326991, 24'd8650311, 24'd8921841, 24'd9087844, 24'd9115470, 24'd8999251, 24'd8762187, 24'd8451192, 24'd8127812, 24'd7856042, 24'd7689667, 24'd7661610, 24'd7777425, 24'd8014192, 24'd8325055, 24'd8648495, 24'd8920503, 24'd9087251, 24'd9115738, 24'd9000328, 24'd8763859, 24'd8453128, 24'd8129629, 24'd7857382, 24'd7690263, 24'd7661345, 24'd7776351, 24'd8012521, 
24'd8323119, 24'd8646676, 24'd8919162, 24'd9086652, 24'd9116001, 24'd9001400, 24'd8765528, 24'd8455064, 24'd8131449, 24'd7858725, 24'd7690864, 24'd7661085, 24'd7775281, 24'd8010854, 24'd8321183, 24'd8644856, 24'd8917817, 24'd9086049, 24'd9116259, 24'd9002467, 24'd8767194, 24'd8457000, 24'd8133270, 24'd7860072, 24'd7691469, 24'd7660829, 24'd7774215, 24'd8009189, 24'd8319248, 24'd8643034, 
24'd8916469, 24'd9085441, 24'd9116511, 24'd9003531, 24'd8768858, 24'd8458934, 24'd8135093, 24'd7861422, 24'd7692080, 24'd7660579, 24'd7773154, 24'd8007526, 24'd8317313, 24'd8641210, 24'd8915116, 24'd9084828, 24'd9116759, 24'd9004590, 24'd8770519, 24'd8460869, 24'd8136918, 24'd7862776, 24'd7692696, 24'd7660334, 24'd7772097, 24'd8005866, 24'd8315379, 24'd8639384, 24'd8913760, 24'd9084210, 
24'd9117001, 24'd9005645, 24'd8772178, 24'd8462803, 24'd8138745, 24'd7864134, 24'd7693316, 24'd7660095, 24'd7771045, 24'd8004209, 24'd8313446, 24'd8637556, 24'd8912400, 24'd9083587, 24'd9117238, 24'd9006695, 24'd8773833, 24'd8464736, 24'd8140573, 24'd7865496, 24'd7693941, 24'd7659860, 24'd7769996, 24'd8002555, 24'd8311512, 24'd8635727, 24'd8911037, 24'd9082959, 24'd9117471, 24'd9007741, 
24'd8775486, 24'd8466669, 24'd8142403, 24'd7866861, 24'd7694571, 24'd7659630, 24'd7768952, 24'd8000903, 24'd8309580, 24'd8633896, 24'd8909670, 24'd9082327, 24'd9117698, 24'd9008783, 24'd8777137, 24'd8468601, 24'd8144235, 24'd7868230, 24'd7695206, 24'd7659406, 24'd7767913, 24'd7999254, 24'd8307648, 24'd8632063, 24'd8908299, 24'd9081689, 24'd9117920, 24'd9009820, 24'd8778784, 24'd8470533, 
24'd8146069, 24'd7869602, 24'd7695846, 24'd7659186, 24'd7766878, 24'd7997608, 24'd8305716, 24'd8630229, 24'd8906925, 24'd9081047, 24'd9118136, 24'd9010853, 24'd8780429, 24'd8472464, 24'd8147904, 24'd7870979, 24'd7696491, 24'd7658972, 24'd7765847, 24'd7995965, 24'd8303786, 24'd8628393, 24'd8905547, 24'd9080400, 24'd9118348, 24'd9011882, 24'd8782071, 24'd8474395, 24'd8149741, 24'd7872358, 
24'd7697141, 24'd7658763, 24'd7764820, 24'd7994324, 24'd8301855, 24'd8626555, 24'd8904165, 24'd9079748, 24'd9118555, 24'd9012906, 24'd8783711, 24'd8476325, 24'd8151579, 24'd7873742, 24'd7697795, 24'd7658559, 24'd7763798, 24'd7992686, 24'd8299926, 24'd8624716, 24'd8902780, 24'd9079091, 24'd9118756, 24'd9013926, 24'd8785347, 24'd8478254, 24'd8153420, 24'd7875129, 24'd7698454, 24'd7658360, 
24'd7762780, 24'd7991051, 24'd8297997, 24'd8622875, 24'd8901391, 24'd9078429, 24'd9118953, 24'd9014942, 24'd8786981, 24'd8480183, 24'd8155262, 24'd7876519, 24'd7699119, 24'd7658166, 24'd7761767, 24'd7989418, 24'd8296068, 24'd8621032, 24'd8899999, 24'd9077763, 24'd9119144, 24'd9015953, 24'd8788612, 24'd8482111, 24'd8157105, 24'd7877914, 24'd7699787, 24'd7657978, 24'd7760758, 24'd7987789, 
24'd8294141, 24'd8619187, 24'd8898603, 24'd9077091, 24'd9119330, 24'd9016960, 24'd8790240, 24'd8484038, 24'd8158950, 24'd7879311, 24'd7700461, 24'd7657794, 24'd7759753, 24'd7986162, 24'd8292213, 24'd8617341, 24'd8897203, 24'd9076415, 24'd9119511, 24'd9017962, 24'd8791866, 24'd8485965, 24'd8160797, 24'd7880713, 24'd7701140, 24'd7657616, 24'd7758753, 24'd7984538, 24'd8290287, 24'd8615494, 
24'd8895800, 24'd9075734, 24'd9119687, 24'd9018960, 24'd8793488, 24'd8487891, 24'd8162646, 24'd7882118, 24'd7701823, 24'd7657442, 24'd7757757, 24'd7982917, 24'd8288361, 24'd8613645, 24'd8894393, 24'd9075048, 24'd9119858, 24'd9019954, 24'd8795108, 24'd8489816, 24'd8164496, 24'd7883526, 24'd7702512, 24'd7657274, 24'd7756766, 24'd7981298, 24'd8286436, 24'd8611794, 24'd8892983, 24'd9074357, 
24'd9120023, 24'd9020943, 24'd8796725, 24'd8491741, 24'd8166347, 24'd7884938, 24'd7703205, 24'd7657111, 24'd7755779, 24'd7979683, 24'd8284512, 24'd8609942, 24'd8891569, 24'd9073662, 24'd9120184, 24'd9021928, 24'd8798339, 24'd8493665, 24'd8168200, 24'd7886354, 24'd7703903, 24'd7656953, 24'd7754797, 24'd7978070, 24'd8282588, 24'd8608088, 24'd8890152, 24'd9072962, 24'd9120339, 24'd9022908, 
24'd8799950, 24'd8495588, 24'd8170055, 24'd7887773, 24'd7704605, 24'd7656800, 24'd7753819, 24'd7976461, 24'd8280666, 24'd8606232, 24'd8888731, 24'd9072257, 24'd9120489, 24'd9023884, 24'd8801558, 24'd8497510, 24'd8171911, 24'd7889195, 24'd7705313, 24'd7656653, 24'd7752845, 24'd7974854, 24'd8278744, 24'd8604375, 24'd8887307, 24'd9071547, 24'd9120634, 24'd9024855, 24'd8803164, 24'd8499432, 
24'd8173769, 24'd7890622, 24'd7706025, 24'd7656510, 24'd7751876, 24'd7973250, 24'd8276822, 24'd8602517, 24'd8885879, 24'd9070832, 24'd9120774, 24'd9025822, 24'd8804766, 24'd8501353, 24'd8175628, 24'd7892051, 24'd7706742, 24'd7656373, 24'd7750911, 24'd7971649, 24'd8274902, 24'd8600657, 24'd8884448, 24'd9070113, 24'd9120909, 24'd9026784, 24'd8806366, 24'd8503273, 24'd8177489, 24'd7893484, 
24'd7707464, 24'd7656240, 24'd7749951, 24'd7970051, 24'd8272982, 24'd8598795, 24'd8883013, 24'd9069389, 24'd9121039, 24'd9027742, 24'd8807962, 24'd8505192, 24'd8179351, 24'd7894921, 24'd7708190, 24'd7656113, 24'd7748995, 24'd7968456, 24'd8271063, 24'd8596932, 24'd8881575, 24'd9068660, 24'd9121163, 24'd9028696, 24'd8809556, 24'd8507111, 24'd8181215, 24'd7896361, 24'd7708922, 24'd7655991, 
24'd7748044, 24'd7966863, 24'd8269145, 24'd8595068, 24'd8880133, 24'd9067926, 24'd9121283, 24'd9029645, 24'd8811147, 24'd8509029, 24'd8183080, 24'd7897804, 24'd7709658, 24'd7655874, 24'd7747098, 24'd7965274, 24'd8267228, 24'd8593202, 24'd8878688, 24'd9067187, 24'd9121397, 24'd9030589, 24'd8812734, 24'd8510945, 24'd8184946, 24'd7899251, 24'd7710399, 24'd7655763, 24'd7746155, 24'd7963688, 
24'd8265311, 24'd8591335, 24'd8877239, 24'd9066444, 24'd9121506, 24'd9031529, 24'd8814319, 24'd8512861, 24'd8186814, 24'd7900701, 24'd7711144, 24'd7655656, 24'd7745218, 24'd7962105, 24'd8263396, 24'd8589466, 24'd8875787, 24'd9065696, 24'd9121610, 24'd9032465, 24'd8815901, 24'd8514776, 24'd8188684, 24'd7902155, 24'd7711895, 24'd7655555, 24'd7744284, 24'd7960524, 24'd8261481, 24'd8587596, 
24'd8874332, 24'd9064943, 24'd9121709, 24'd9033396, 24'd8817480, 24'd8516691, 24'd8190554, 24'd7903612, 24'd7712650, 24'd7655458, 24'd7743356, 24'd7958947, 24'd8259568, 24'd8585725, 24'd8872873, 24'd9064186, 24'd9121803, 24'd9034322, 24'd8819055, 24'd8518604, 24'd8192427, 24'd7905073, 24'd7713410, 24'd7655367, 24'd7742431, 24'd7957373, 24'd8257655, 24'd8583852, 24'd8871411, 24'd9063423, 
24'd9121891, 24'd9035244, 24'd8820628, 24'd8520516, 24'd8194300, 24'd7906537, 24'd7714174, 24'd7655281, 24'd7741512, 24'd7955802, 24'd8255743, 24'd8581978, 24'd8869945, 24'd9062656, 24'd9121975, 24'd9036161, 24'd8822198, 24'd8522428, 24'd8196175, 24'd7908004, 24'd7714944, 24'd7655200, 24'd7740597, 24'd7954233, 24'd8253832, 24'd8580102, 24'd8868476, 24'd9061885, 24'd9122053, 24'd9037074, 
24'd8823765, 24'd8524338, 24'd8198051, 24'd7909475, 24'd7715718, 24'd7655125, 24'd7739686, 24'd7952668, 24'd8251922, 24'd8578225, 24'd8867004, 24'd9061108, 24'd9122126, 24'd9037982, 24'd8825328, 24'd8526248, 24'd8199929, 24'd7910949, 24'd7716497, 24'd7655054, 24'd7738780, 24'd7951106, 24'd8250013, 24'd8576347, 24'd8865528, 24'd9060327, 24'd9122194, 24'd9038886, 24'd8826889, 24'd8528157, 
24'd8201808, 24'd7912426, 24'd7717280, 24'd7654989, 24'd7737879, 24'd7949547, 24'd8248104, 24'd8574467, 24'd8864049, 24'd9059541, 24'd9122257, 24'd9039785, 24'd8828446, 24'd8530064, 24'd8203688, 24'd7913907, 24'd7718068, 24'd7654928, 24'd7736982, 24'd7947991, 24'd8246197, 24'd8572586, 24'd8862566, 24'd9058751, 24'd9122315, 24'd9040680, 24'd8830001, 24'd8531971, 24'd8205570, 24'd7915391, 
24'd7718861, 24'd7654873, 24'd7736090, 24'd7946438, 24'd8244291, 24'd8570704, 24'd8861081, 24'd9057955, 24'd9122368, 24'd9041570, 24'd8831552, 24'd8533877, 24'd8207452, 24'd7916878, 24'd7719659, 24'd7654823, 24'd7735202, 24'd7944888, 24'd8242386, 24'd8568821, 24'd8859592, 24'd9057156, 24'd9122415, 24'd9042455, 24'd8833100, 24'd8535781, 24'd8209336, 24'd7918369, 24'd7720461, 24'd7654778, 
24'd7734319, 24'd7943342, 24'd8240482, 24'd8566936, 24'd8858099, 24'd9056351, 24'd9122457, 24'd9043336, 24'd8834646, 24'd8537685, 24'd8211222, 24'd7919863, 24'd7721268, 24'd7654738, 24'd7733440, 24'd7941798, 24'd8238579, 24'd8565050, 24'd8856604, 24'd9055542, 24'd9122494, 24'd9044213, 24'd8836188, 24'd8539587, 24'd8213108, 24'd7921360, 24'd7722080, 24'd7654704, 24'd7732566, 24'd7940258, 
24'd8236677, 24'd8563163, 24'd8855105, 24'd9054728, 24'd9122527, 24'd9045084, 24'd8837726, 24'd8541489, 24'd8214996, 24'd7922861, 24'd7722896, 24'd7654674, 24'd7731697, 24'd7938720, 24'd8234776, 24'd8561274, 24'd8853602, 24'd9053909, 24'd9122553, 24'd9045951, 24'd8839262, 24'd8543389, 24'd8216885, 24'd7924365, 24'd7723717, 24'd7654650, 24'd7730832, 24'd7937186, 24'd8232876, 24'd8559385, 
24'd8852097, 24'd9053086, 24'd9122575, 24'd9046814, 24'd8840795, 24'd8545289, 24'd8218775, 24'd7925872, 24'd7724543, 24'd7654631, 24'd7729972, 24'd7935655, 24'd8230977, 24'd8557494, 24'd8850588, 24'd9052258, 24'd9122592, 24'd9047672, 24'd8842324, 24'd8547187, 24'd8220667, 24'd7927382, 24'd7725373, 24'd7654617, 24'd7729116, 24'd7934127, 24'd8229080, 24'd8555602, 24'd8849076, 24'd9051425, 
24'd9122603, 24'd9048525, 24'd8843850, 24'd8549084, 24'd8222560, 24'd7928896, 24'd7726208, 24'd7654608, 24'd7728265, 24'd7932603, 24'd8227183, 24'd8553709, 24'd8847561, 24'd9050588, 24'd9122609, 24'd9049373, 24'd8845373, 24'd8550980, 24'd8224453, 24'd7930413, 24'd7727048, 24'd7654604, 24'd7727419, 24'd7931081, 24'd8225288, 24'd8551814, 24'd8846043, 24'd9049746, 24'd9122610, 24'd9050217, 
24'd8846893, 24'd8552875, 24'd8226348, 24'd7931933, 24'd7727892, 24'd7654606, 24'd7726577, 24'd7929563, 24'd8223393, 24'd8549919, 24'd8844521, 24'd9048899, 24'd9122606, 24'd9051057, 24'd8848410, 24'd8554768, 24'd8228244, 24'd7933456, 24'd7728741, 24'd7654612, 24'd7725740, 24'd7928048, 24'd8221500, 24'd8548022, 24'd8842996, 24'd9048048, 24'd9122597, 24'd9051891, 24'd8849923, 24'd8556661, 
24'd8230141, 24'd7934982, 24'd7729594, 24'd7654624, 24'd7724908, 24'd7926537, 24'd8219608, 24'd8546125, 24'd8841468, 24'd9047192, 24'd9122583, 24'd9052722, 24'd8851433, 24'd8558552, 24'd8232040, 24'd7936512, 24'd7730453, 24'd7654641, 24'd7724080, 24'd7925028, 24'd8217717, 24'd8544226, 24'd8839937, 24'd9046332, 24'd9122564, 24'd9053547, 24'd8852940, 24'd8560442, 24'd8233939, 24'd7938044, 
24'd7731315, 24'd7654663, 24'd7723257, 24'd7923523, 24'd8215828, 24'd8542326, 24'd8838403, 24'd9045467, 24'd9122539, 24'd9054368, 24'd8854444, 24'd8562331, 24'd8235840, 24'd7939580, 24'd7732183, 24'd7654690, 24'd7722439, 24'd7922021, 24'd8213940, 24'd8540425, 24'd8836866, 24'd9044597, 24'd9122509, 24'd9055184, 24'd8855944, 24'd8564219, 24'd8237741, 24'd7941119, 24'd7733055, 24'd7654723, 
24'd7721625, 24'd7920522, 24'd8212052, 24'd8538523, 24'd8835325, 24'd9043723, 24'd9122474, 24'd9055995, 24'd8857441, 24'd8566106, 24'd8239644, 24'd7942662, 24'd7733931, 24'd7654760, 24'd7720816, 24'd7919027, 24'd8210167, 24'd8536620, 24'd8833781, 24'd9042844, 24'd9122434, 24'd9056802, 24'd8858935, 24'd8567991, 24'd8241547, 24'd7944207, 24'd7734812, 24'd7654803, 24'd7720012, 24'd7917535, 
24'd8208282, 24'd8534715, 24'd8832234, 24'd9041960, 24'd9122389, 24'd9057604, 24'd8860425, 24'd8569875, 24'd8243452, 24'd7945755, 24'd7735698, 24'd7654850, 24'd7719212, 24'd7916046, 24'd8206399, 24'd8532810, 24'd8830684, 24'd9041072, 24'd9122339, 24'd9058401, 24'd8861913, 24'd8571758, 24'd8245358, 24'd7947307, 24'd7736588, 24'd7654903, 24'd7718417, 24'd7914560, 24'd8204516, 24'd8530904, 
24'd8829131, 24'd9040180, 24'd9122283, 24'd9059194, 24'd8863396, 24'd8573639, 24'd8247265, 24'd7948861, 24'd7737483, 24'd7654961, 24'd7717627, 24'd7913078, 24'd8202636, 24'd8528997, 24'd8827575, 24'd9039283, 24'd9122223, 24'd9059982, 24'd8864877, 24'd8575519, 24'd8249172, 24'd7950419, 24'd7738383, 24'd7655025, 24'd7716841, 24'd7911599, 24'd8200756, 24'd8527089, 24'd8826016, 24'd9038381, 
24'd9122157, 24'd9060765, 24'd8866354, 24'd8577398, 24'd8251081, 24'd7951980, 24'd7739287, 24'd7655093, 24'd7716060, 24'd7910124, 24'd8198878, 24'd8525179, 24'd8824454, 24'd9037475, 24'd9122086, 24'd9061543, 24'd8867828, 24'd8579276, 24'd8252991, 24'd7953544, 24'd7740195, 24'd7655166, 24'd7715284, 24'd7908651, 24'd8197001, 24'd8523269, 24'd8822888, 24'd9036564, 24'd9122010, 24'd9062317, 
24'd8869298, 24'd8581152, 24'd8254901, 24'd7955111, 24'd7741108, 24'd7655245, 24'd7714513, 24'd7907183, 24'd8195126, 24'd8521358, 24'd8821320, 24'd9035648, 24'd9121929, 24'd9063086, 24'd8870766, 24'd8583027, 24'd8256813, 24'd7956681, 24'd7742026, 24'd7655329, 24'd7713746, 24'd7905717, 24'd8193251, 24'd8519446, 24'd8819748, 24'd9034729, 24'd9121842, 24'd9063851, 24'd8872229, 24'd8584900, 
24'd8258725, 24'd7958253, 24'd7742948, 24'd7655418, 24'd7712984, 24'd7904255, 24'd8191379, 24'd8517533, 24'd8818174, 24'd9033804, 24'd9121751, 24'd9064610, 24'd8873690, 24'd8586772, 24'd8260638, 24'd7959829, 24'd7743875, 24'd7655512, 24'd7712227, 24'd7902796, 24'd8189507, 24'd8515620, 24'd8816596, 24'd9032875, 24'd9121654, 24'd9065365, 24'd8875147, 24'd8588643, 24'd8262553, 24'd7961408, 
24'd7744806, 24'd7655611, 24'd7711474, 24'd7901341, 24'd8187637, 24'd8513705, 24'd8815016, 24'd9031942, 24'd9121553, 24'd9066115, 24'd8876600, 24'd8590512, 24'd8264468, 24'd7962990, 24'd7745742, 24'd7655715, 24'd7710727, 24'd7899889, 24'd8185769, 24'd8511789, 24'd8813432, 24'd9031004, 24'd9121446, 24'd9066861, 24'd8878050, 24'd8592380, 24'd8266384, 24'd7964575, 24'd7746682, 24'd7655825, 
24'd7709984, 24'd7898441, 24'd8183901, 24'd8509873, 24'd8811846, 24'd9030061, 24'd9121334, 24'd9067601, 24'd8879497, 24'd8594247, 24'd8268301, 24'd7966163, 24'd7747627, 24'd7655939, 24'd7709245, 24'd7896996, 24'd8182036, 24'd8507956, 24'd8810257, 24'd9029114, 24'd9121217, 24'd9068337, 24'd8880940, 24'd8596112, 24'd8270218, 24'd7967754, 24'd7748576, 24'd7656059, 24'd7708512, 24'd7895554, 
24'd8180171, 24'd8506037, 24'd8808664, 24'd9028163, 24'd9121094, 24'd9069068, 24'd8882380, 24'd8597975, 24'd8272137, 24'd7969348, 24'd7749530, 24'd7656184, 24'd7707783, 24'd7894116, 24'd8178309, 24'd8504118, 24'd8807069, 24'd9027207, 24'd9120967, 24'd9069794, 24'd8883816, 24'd8599837, 24'd8274056, 24'd7970945, 24'd7750488, 24'd7656314, 24'd7707059, 24'd7892682, 24'd8176447, 24'd8502199, 
24'd8805471, 24'd9026246, 24'd9120834, 24'd9070516, 24'd8885249, 24'd8601698, 24'd8275977, 24'd7972545, 24'd7751451, 24'd7656449, 24'd7706340, 24'd7891251, 24'd8174587, 24'd8500278, 24'd8803870, 24'd9025281, 24'd9120697, 24'd9071233, 24'd8886679, 24'd8603557, 24'd8277897, 24'd7974147, 24'd7752418, 24'd7656589, 24'd7705626, 24'd7889823, 24'd8172729, 24'd8498357, 24'd8802265, 24'd9024312, 
24'd9120554, 24'd9071945, 24'd8888104, 24'd8605415, 24'd8279819, 24'd7975753, 24'd7753389, 24'd7656735, 24'd7704916, 24'd7888399, 24'd8170872, 24'd8496435, 24'd8800658, 24'd9023338, 24'd9120406, 24'd9072652, 24'd8889527, 24'd8607271, 24'd8281742, 24'd7977361, 24'd7754365, 24'd7656885, 24'd7704211, 24'd7886978, 24'd8169017, 24'd8494512, 24'd8799049, 24'd9022360, 24'd9120253, 24'd9073354, 
24'd8890946, 24'd8609125, 24'd8283665, 24'd7978972, 24'd7755346, 24'd7657041, 24'd7703511, 24'd7885561, 24'd8167163, 24'd8492588, 24'd8797436, 24'd9021377, 24'd9120094, 24'd9074052, 24'd8892361, 24'd8610978, 24'd8285589, 24'd7980587, 24'd7756331, 24'd7657202, 24'd7702816, 24'd7884148, 24'd8165311, 24'd8490664, 24'd8795820, 24'd9020390, 24'd9119931, 24'd9074745, 24'd8893773, 24'd8612830, 
24'd8287514, 24'd7982204, 24'd7757320, 24'd7657368, 24'd7702126, 24'd7882738, 24'd8163460, 24'd8488739, 24'd8794202, 24'd9019398, 24'd9119763, 24'd9075433, 24'd8895181, 24'd8614680, 24'd8289439, 24'd7983824, 24'd7758314, 24'd7657539, 24'd7701440, 24'd7881331, 24'd8161611, 24'd8486813, 24'd8792580, 24'd9018402, 24'd9119589, 24'd9076116, 24'd8896586, 24'd8616528, 24'd8291365, 24'd7985446, 
24'd7759312, 24'd7657715, 24'd7700759, 24'd7879928, 24'd8159763, 24'd8484887, 24'd8790956, 24'd9017402, 24'd9119410, 24'd9076794, 24'd8897987, 24'd8618375, 24'd8293292, 24'd7987072, 24'd7760315, 24'd7657896, 24'd7700084, 24'd7878529, 24'd8157918, 24'd8482959, 24'd8789329, 24'd9016397, 24'd9119226, 24'd9077468, 24'd8899385, 24'd8620220, 24'd8295219, 24'd7988700, 24'd7761322, 24'd7658082, 
24'd7699412, 24'd7877133, 24'd8156073, 24'd8481032, 24'd8787700, 24'd9015388, 24'd9119037, 24'd9078136, 24'd8900779, 24'd8622063, 24'd8297147, 24'd7990331, 24'd7762333, 24'd7658274, 24'd7698746, 24'd7875741, 24'd8154231, 24'd8479103, 24'd8786067, 24'd9014374, 24'd9118843, 24'd9078800, 24'd8902169, 24'd8623905, 24'd8299076, 24'd7991965, 24'd7763349, 24'd7658471, 24'd7698085, 24'd7874352, 
24'd8152390, 24'd8477174, 24'd8784432, 24'd9013356, 24'd9118644, 24'd9079459, 24'd8903556, 24'd8625745, 24'd8301006, 24'd7993602, 24'd7764370, 24'd7658672, 24'd7697428, 24'd7872967, 24'd8150550, 24'd8475245, 24'd8782793, 24'd9012334, 24'd9118440, 24'd9080113, 24'd8904939, 24'd8627584, 24'd8302936, 24'd7995242, 24'd7765394, 24'd7658879, 24'd7696776, 24'd7871586, 24'd8148713, 24'd8473314, 
24'd8781153, 24'd9011307, 24'd9118230, 24'd9080763, 24'd8906319, 24'd8629421, 24'd8304866, 24'd7996884, 24'd7766423, 24'd7659091, 24'd7696130, 24'd7870208, 24'd8146877, 24'd8471383, 24'd8779509, 24'd9010276, 24'd9118016, 24'd9081407, 24'd8907695, 24'd8631256, 24'd8306797, 24'd7998529, 24'd7767456, 24'd7659309, 24'd7695488, 24'd7868834, 24'd8145042, 24'd8469452, 24'd8777862, 24'd9009240, 
24'd9117796, 24'd9082047, 24'd8909067, 24'd8633089, 24'd8308729, 24'd8000177, 24'd7768494, 24'd7659531, 24'd7694850, 24'd7867463, 24'd8143210, 24'd8467520, 24'd8776213, 24'd9008200, 24'd9117571, 24'd9082681, 24'd8910436, 24'd8634921, 24'd8310661, 24'd8001827, 24'd7769536, 24'd7659758, 24'd7694218, 24'd7866096, 24'd8141379, 24'd8465587, 24'd8774562, 24'd9007156, 24'd9117341, 24'd9083311, 
24'd8911801, 24'd8636751, 24'd8312594, 24'd8003480, 24'd7770583, 24'd7659991, 24'd7693591, 24'd7864733, 24'd8139550, 24'd8463654, 24'd8772907, 24'd9006108, 24'd9117106, 24'd9083936, 24'd8913162, 24'd8638579, 24'd8314528, 24'd8005136, 24'd7771633, 24'd7660228, 24'd7692968, 24'd7863374, 24'd8137722, 24'd8461720, 24'd8771250, 24'd9005055, 24'd9116866, 24'd9084556, 24'd8914520, 24'd8640406, 
24'd8316462, 24'd8006795, 24'd7772688, 24'd7660471, 24'd7692350, 24'd7862018, 24'd8135897, 24'd8459786, 24'd8769590, 24'd9003998, 24'd9116621, 24'd9085172, 24'd8915874, 24'd8642231, 24'd8318396, 24'd8008456, 24'd7773748, 24'd7660719, 24'd7691738, 24'd7860666, 24'd8134073, 24'd8457852, 24'd8767927, 24'd9002936, 24'd9116371, 24'd9085782, 24'd8917224, 24'd8644054, 24'd8320331, 24'd8010120, 
24'd7774811, 24'd7660972, 24'd7691130, 24'd7859317, 24'd8132251, 24'd8455916, 24'd8766262, 24'd9001870, 24'd9116115, 24'd9086387, 24'd8918570, 24'd8645875, 24'd8322266, 24'd8011787, 24'd7775879, 24'd7661230, 24'd7690527, 24'd7857973, 24'd8130430, 24'd8453981, 24'd8764594, 24'd9000800, 24'd9115855, 24'd9086988, 24'd8919913, 24'd8647694, 24'd8324202, 24'd8013456, 24'd7776951, 24'd7661493, 
24'd7689929, 24'd7856632, 24'd8128612, 24'd8452045, 24'd8762923, 24'd8999726, 24'd9115589, 24'd9087584, 24'd8921252, 24'd8649512, 24'd8326138, 24'd8015128, 24'd7778028, 24'd7661761, 24'd7689335, 24'd7855294, 24'd8126795, 24'd8450108, 24'd8761250, 24'd8998647, 24'd9115318, 24'd9088174, 24'd8922588, 24'd8651327, 24'd8328075, 24'd8016802, 24'd7779109, 24'd7662034, 24'd7688747, 24'd7853961, 
24'd8124980, 24'd8448171, 24'd8759575, 24'd8997564, 24'd9115042, 24'd9088760, 24'd8923919, 24'd8653141, 24'd8330012, 24'd8018479, 24'd7780194, 24'd7662313, 24'd7688164, 24'd7852631, 24'd8123167, 24'd8446234, 24'd8757896, 24'd8996477, 24'd9114761, 24'd9089341, 24'd8925247, 24'd8654953, 24'd8331950, 24'd8020159, 24'd7781283, 24'd7662596, 24'd7687585, 24'd7851305, 24'd8121356, 24'd8444296, 
24'd8756215, 24'd8995385, 24'd9114475, 24'd9089917, 24'd8926571, 24'd8656763, 24'd8333888, 24'd8021841, 24'd7782377, 24'd7662885, 24'd7687011, 24'd7849983, 24'd8119547, 24'd8442358, 24'd8754532, 24'd8994290, 24'd9114184, 24'd9090488, 24'd8927892, 24'd8658572, 24'd8335826, 24'd8023526, 24'd7783475, 24'd7663178, 24'd7686443, 24'd7848664, 24'd8117740, 24'd8440419, 24'd8752846, 24'd8993190, 
24'd9113888, 24'd9091055, 24'd8929208, 24'd8660378, 24'd8337765, 24'd8025213, 24'd7784577, 24'd7663477, 24'd7685879, 24'd7847350, 24'd8115934, 24'd8438481, 24'd8751157, 24'd8992085, 24'd9113587, 24'd9091616, 24'd8930521, 24'd8662183, 24'd8339704, 24'd8026903, 24'd7785683, 24'd7663781, 24'd7685320, 24'd7846039, 24'd8114131, 24'd8436541, 24'd8749466, 24'd8990977, 24'd9113280, 24'd9092172, 
24'd8931830, 24'd8663985, 24'd8341644, 24'd8028596, 24'd7786794, 24'd7664090, 24'd7684766, 24'd7844732, 24'd8112329, 24'd8434602, 24'd8747772, 24'd8989864, 24'd9112969, 24'd9092724, 24'd8933135, 24'd8665786, 24'd8343583, 24'd8030291, 24'd7787909, 24'd7664404, 24'd7684217, 24'd7843428, 24'd8110530, 24'd8432662, 24'd8746076, 24'd8988747, 24'd9112652, 24'd9093270, 24'd8934437, 24'd8667585, 
24'd8345523, 24'd8031988, 24'd7789028, 24'd7664723, 24'd7683673, 24'd7842129, 24'd8108732, 24'd8430722, 24'd8744377, 24'd8987626, 24'd9112331, 24'd9093812, 24'd8935734, 24'd8669381, 24'd8347464, 24'd8033688, 24'd7790151, 24'd7665047, 24'd7683134, 24'd7840833, 24'd8106936, 24'd8428781, 24'd8742676, 24'd8986501, 24'd9112004, 24'd9094348, 24'd8937028, 24'd8671176, 24'd8349404, 24'd8035391, 
24'd7791278, 24'd7665376, 24'd7682600, 24'd7839542, 24'd8105142, 24'd8426840, 24'd8740972, 24'd8985371, 24'd9111672, 24'd9094880, 24'd8938318, 24'd8672969, 24'd8351345, 24'd8037096, 24'd7792410, 24'd7665710, 24'd7682071, 24'd7838254, 24'd8103350, 24'd8424899, 24'd8739266, 24'd8984238, 24'd9111336, 24'd9095407, 24'd8939604, 24'd8674760, 24'd8353287, 24'd8038803, 24'd7793546, 24'd7666050, 
24'd7681547, 24'd7836970, 24'd8101561, 24'd8422958, 24'd8737557, 24'd8983100, 24'd9110994, 24'd9095929, 24'd8940886, 24'd8676548, 24'd8355228, 24'd8040513, 24'd7794686, 24'd7666394, 24'd7681027, 24'd7835689, 24'd8099773, 24'd8421016, 24'd8735846, 24'd8981958, 24'd9110647, 24'd9096445, 24'd8942164, 24'd8678335, 24'd8357170, 24'd8042226, 24'd7795830, 24'd7666744, 24'd7680513, 24'd7834413, 
24'd8097987, 24'd8419074, 24'd8734132, 24'd8980812, 24'd9110295, 24'd9096957, 24'd8943439, 24'd8680120, 24'd8359112, 24'd8043940, 24'd7796978, 24'd7667098, 24'd7680004, 24'd7833141, 24'd8096203, 24'd8417132, 24'd8732416, 24'd8979661, 24'd9109938, 24'd9097464, 24'd8944709, 24'd8681903, 24'd8361054, 24'd8045657, 24'd7798131, 24'd7667458, 24'd7679499, 24'd7831872, 24'd8094422, 24'd8415190, 
24'd8730698, 24'd8978507, 24'd9109575, 24'd9097966, 24'd8945976, 24'd8683683, 24'd8362996, 24'd8047377, 24'd7799287, 24'd7667823, 24'd7679000, 24'd7830607, 24'd8092642, 24'd8413248, 24'd8728977, 24'd8977348, 24'd9109208, 24'd9098463, 24'd8947238, 24'd8685462, 24'd8364938, 24'd8049099, 24'd7800448, 24'd7668192, 24'd7678506, 24'd7829347, 24'd8090865, 24'd8411305, 24'd8727254, 24'd8976185, 
24'd9108836, 24'd9098955, 24'd8948497, 24'd8687238, 24'd8366881, 24'd8050823, 24'd7801613, 24'd7668567, 24'd7678016, 24'd7828090, 24'd8089089, 24'd8409363, 24'd8725529, 24'd8975018, 24'd9108459, 24'd9099442, 24'd8949752, 24'd8689013, 24'd8368824, 24'd8052550, 24'd7802782, 24'd7668947, 24'd7677532, 24'd7826837, 24'd8087316, 24'd8407420, 24'd8723801, 24'd8973847, 24'd9108076, 24'd9099924, 
24'd8951003, 24'd8690785, 24'd8370767, 24'd8054279, 24'd7803955, 24'd7669332, 24'd7677052, 24'd7825588, 24'd8085545, 24'd8405477, 24'd8722070, 24'd8972672, 24'd9107689, 24'd9100401, 24'd8952250, 24'd8692555, 24'd8372710, 24'd8056011, 24'd7805132, 24'd7669722, 24'd7676578, 24'd7824343, 24'd8083775, 24'd8403534, 24'd8720338, 24'd8971493, 24'd9107297, 24'd9100873, 24'd8953493, 24'd8694323, 
24'd8374653, 24'd8057744, 24'd7806313, 24'd7670117, 24'd7676108, 24'd7823102, 24'd8082009, 24'd8401590, 24'd8718603, 24'd8970310, 24'd9106899, 24'd9101340, 24'd8954732, 24'd8696089, 24'd8376596, 24'd8059480, 24'd7807498, 24'd7670517, 24'd7675644, 24'd7821865, 24'd8080244, 24'd8399647, 24'd8716866, 24'd8969123, 24'd9106497, 24'd9101802, 24'd8955967, 24'd8697853, 24'd8378540, 24'd8061219, 
24'd7808688, 24'd7670922, 24'd7675184, 24'd7820632, 24'd8078481, 24'd8397704, 24'd8715126, 24'd8967931, 24'd9106089, 24'd9102259, 24'd8957198, 24'd8699614, 24'd8380483, 24'd8062960, 24'd7809881, 24'd7671332, 24'd7674730, 24'd7819403, 24'd8076721, 24'd8395760, 24'd8713384, 24'd8966736, 24'd9105677, 24'd9102711, 24'd8958425, 24'd8701374, 24'd8382427, 24'd8064703, 24'd7811079, 24'd7671747, 
24'd7674280, 24'd7818178, 24'd8074962, 24'd8393817, 24'd8711640, 24'd8965536, 24'd9105259, 24'd9103158, 24'd8959648, 24'd8703131, 24'd8384370, 24'd8066448, 24'd7812280, 24'd7672167, 24'd7673836, 24'd7816957, 24'd8073206, 24'd8391873, 24'd8709894, 24'd8964333, 24'd9104836, 24'd9103600, 24'd8960868, 24'd8704886, 24'd8386314, 24'd8068195, 24'd7813486, 24'd7672592, 24'd7673396, 24'd7815739, 
24'd8071452, 24'd8389930, 24'd8708145, 24'd8963125, 24'd9104409, 24'd9104037, 24'd8962083, 24'd8706639, 24'd8388257, 24'd8069945, 24'd7814695, 24'd7673022, 24'd7672962, 24'd7814526, 24'd8069701, 24'd8387986, 24'd8706394, 24'd8961913, 24'd9103976, 24'd9104469, 24'd8963294, 24'd8708389, 24'd8390201, 24'd8071697, 24'd7815909, 24'd7673457, 24'd7672532, 24'd7813317, 24'd8067951, 24'd8386042, 
24'd8704641, 24'd8960698, 24'd9103538, 24'd9104896, 24'd8964501, 24'd8710138, 24'd8392144, 24'd8073451, 24'd7817127, 24'd7673897, 24'd7672108, 24'd7812112, 24'd8066204, 24'd8384099, 24'd8702886, 24'd8959478, 24'd9103096, 24'd9105318, 24'd8965704, 24'd8711884, 24'd8394088, 24'd8075208, 24'd7818348, 24'd7674343, 24'd7671688, 24'd7810911, 24'd8064459, 24'd8382155, 24'd8701128, 24'd8958254, 
24'd9102648, 24'd9105734, 24'd8966903, 24'd8713628, 24'd8396031, 24'd8076966, 24'd7819574, 24'd7674793, 24'd7671274, 24'd7809714, 24'd8062716, 24'd8380212, 24'd8699369, 24'd8957027, 24'd9102195, 24'd9106146, 24'd8968098, 24'd8715369, 24'd8397975, 24'd8078727, 24'd7820804, 24'd7675248, 24'd7670865, 24'd7808521, 24'd8060976, 24'd8378268, 24'd8697607, 24'd8955795, 24'd9101738, 24'd9106553, 
24'd8969289, 24'd8717108, 24'd8399918, 24'd8080490, 24'd7822037, 24'd7675708, 24'd7670460, 24'd7807333, 24'd8059238, 24'd8376325, 24'd8695843, 24'd8954559, 24'd9101275, 24'd9106955, 24'd8970475, 24'd8718845, 24'd8401862, 24'd8082255, 24'd7823275, 24'd7676173, 24'd7670061, 24'd7806148, 24'd8057502, 24'd8374382, 24'd8694077, 24'd8953320, 24'd9100807, 24'd9107352, 24'd8971658, 24'd8720580, 
24'd8403805, 24'd8084022, 24'd7824517, 24'd7676644, 24'd7669667, 24'd7804967, 24'd8055769, 24'd8372439, 24'd8692308, 24'd8952076, 24'd9100334, 24'd9107743, 24'd8972837, 24'd8722312, 24'd8405748, 24'd8085792, 24'd7825762, 24'd7677119, 24'd7669278, 24'd7803791, 24'd8054038, 24'd8370496, 24'd8690538, 24'd8950829, 24'd9099857, 24'd9108130, 24'd8974011, 24'd8724042, 24'd8407691, 24'd8087563, 
24'd7827012, 24'd7677599, 24'd7668893, 24'd7802618, 24'd8052309, 24'd8368553, 24'd8688765, 24'd8949577, 24'd9099374, 24'd9108512, 24'd8975182, 24'd8725770, 24'd8409634, 24'd8089337, 24'd7828265, 24'd7678084, 24'd7668514, 24'd7801450, 24'd8050583, 24'd8366610, 24'd8686991, 24'd8948322, 24'd9098886, 24'd9108888, 24'd8976348, 24'd8727495, 24'd8411576, 24'd8091113, 24'd7829523, 24'd7678574, 
24'd7668140, 24'd7800285, 24'd8048859, 24'd8364667, 24'd8685214, 24'd8947062, 24'd9098394, 24'd9109260, 24'd8977510, 24'd8729218, 24'd8413519, 24'd8092890, 24'd7830784, 24'd7679069, 24'd7667771, 24'd7799125, 24'd8047137, 24'd8362725, 24'd8683435, 24'd8945799, 24'd9097896, 24'd9109626, 24'd8978668, 24'd8730938, 24'd8415461, 24'd8094670, 24'd7832049, 24'd7679569, 24'd7667407, 24'd7797969, 
24'd8045418, 24'd8360783, 24'd8681654, 24'd8944532, 24'd9097394, 24'd9109988, 24'd8979822, 24'd8732656, 24'd8417404, 24'd8096452, 24'd7833318, 24'd7680075, 24'd7667048, 24'd7796818, 24'd8043701, 24'd8358840, 24'd8679871, 24'd8943261, 24'd9096886, 24'd9110344, 24'd8980972, 24'd8734372, 24'd8419346, 24'd8098236, 24'd7834591, 24'd7680585, 24'd7666695, 24'd7795670, 24'd8041986, 24'd8356899, 
24'd8678086, 24'd8941986, 24'd9096374, 24'd9110695, 24'd8982117, 24'd8736085, 24'd8421287, 24'd8100022, 24'd7835868, 24'd7681100, 24'd7666346, 24'd7794526, 24'd8040274, 24'd8354957, 24'd8676299, 24'd8940707, 24'd9095856, 24'd9111042, 24'd8983259, 24'd8737796, 24'd8423229, 24'd8101810, 24'd7837149, 24'd7681620, 24'd7666002, 24'd7793387, 24'd8038565, 24'd8353016, 24'd8674510, 24'd8939425, 
24'd9095334, 24'd9111383, 24'd8984396, 24'd8739504, 24'd8425170, 24'd8103601, 24'd7838433, 24'd7682144, 24'd7665663, 24'd7792252, 24'd8036858, 24'd8351074, 24'd8672719, 24'd8938138, 24'd9094806, 24'd9111719, 24'd8985529, 24'd8741210, 24'd8427111, 24'd8105393, 24'd7839722, 24'd7682674, 24'd7665330, 24'd7791121, 24'd8035153, 24'd8349133, 24'd8670926, 24'd8936848, 24'd9094274, 24'd9112050, 
24'd8986658, 24'd8742913, 24'd8429052, 24'd8107187, 24'd7841014, 24'd7683209, 24'd7665001, 24'd7789994, 24'd8033451, 24'd8347193, 24'd8669131, 24'd8935553, 24'd9093737, 24'd9112376, 24'd8987783, 24'd8744614, 24'd8430992, 24'd8108983, 24'd7842310, 24'd7683749, 24'd7664678, 24'd7788871, 24'd8031751, 24'd8345252, 24'd8667334, 24'd8934255, 24'd9093194, 24'd9112697, 24'd8988903, 24'd8746313, 
24'd8432933, 24'd8110781, 24'd7843610, 24'd7684294, 24'd7664360, 24'd7787753, 24'd8030054, 24'd8343312, 24'd8665535, 24'd8932953, 24'd9092647, 24'd9113013, 24'd8990020, 24'd8748009, 24'd8434872, 24'd8112581, 24'd7844914, 24'd7684843, 24'd7664046, 24'd7786639, 24'd8028359, 24'd8341373, 24'd8663734, 24'd8931648, 24'd9092095, 24'd9113323, 24'd8991132, 24'd8749702, 24'd8436812, 24'd8114382, 
24'd7846222, 24'd7685398, 24'd7663738, 24'd7785529, 24'd8026667, 24'd8339433, 24'd8661931, 24'd8930338, 24'd9091538, 24'd9113629, 24'd8992240, 24'd8751393, 24'd8438751, 24'd8116186, 24'd7847533, 24'd7685957, 24'd7663435, 24'd7784423, 24'd8024978, 24'd8337494, 24'd8660126, 24'd8929025, 24'd9090976, 24'd9113930, 24'd8993343, 24'd8753081, 24'd8440690, 24'd8117992, 24'd7848848, 24'd7686522, 
24'd7663137, 24'd7783321, 24'd8023291, 24'd8335556, 24'd8658319, 24'd8927708, 24'd9090409, 24'd9114225, 24'd8994443, 24'd8754767, 24'd8442629, 24'd8119800, 24'd7850167, 24'd7687091, 24'd7662844, 24'd7782224, 24'd8021606, 24'd8333617, 24'd8656511, 24'd8926387, 24'd9089837, 24'd9114516, 24'd8995538, 24'd8756450, 24'd8444567, 24'd8121609, 24'd7851490, 24'd7687666, 24'd7662556, 24'd7781131, 
24'd8019924, 24'd8331679, 24'd8654700, 24'd8925062, 24'd9089260, 24'd9114801, 24'd8996629, 24'd8758131, 24'd8446504, 24'd8123420, 24'd7852817, 24'd7688245, 24'd7662273, 24'd7780042, 24'd8018245, 24'd8329742, 24'd8652888, 24'd8923734, 24'd9088679, 24'd9115081, 24'd8997716, 24'd8759809, 24'd8448442, 24'd8125234, 24'd7854147, 24'd7688829, 24'd7661996, 24'd7778958, 24'd8016568, 24'd8327805, 
24'd8651074, 24'd8922402, 24'd9088092, 24'd9115356, 24'd8998798, 24'd8761484, 24'd8450379, 24'd8127049, 24'd7855481, 24'd7689418, 24'd7661723, 24'd7777877, 24'd8014894, 24'd8325868, 24'd8649258, 24'd8921066, 24'd9087501, 24'd9115626, 24'd8999876, 24'd8763157, 24'd8452315, 24'd8128866, 24'd7856819, 24'd7690012, 24'd7661456, 24'd7776802, 24'd8013223, 24'd8323932, 24'd8647440, 24'd8919726, 
24'd9086904, 24'd9115891, 24'd9000950, 24'd8764827, 24'd8454251, 24'd8130684, 24'd7858160, 24'd7690611, 24'd7661193, 24'd7775730, 24'd8011554, 24'd8321996, 24'd8645621, 24'd8918383, 24'd9086303, 24'd9116151, 24'd9002019, 24'd8766495, 24'd8456187, 24'd8132505, 24'd7859505, 24'd7691214, 24'd7660936, 24'd7774663, 24'd8009888, 24'd8320061, 24'd8643799, 24'd8917036, 24'd9085697, 24'd9116406, 
24'd9003085, 24'd8768159, 24'd8458122, 24'd8134327, 24'd7860854, 24'd7691823, 24'd7660684, 24'd7773599, 24'd8008224, 24'd8318126, 24'd8641976, 24'd8915685, 24'd9085086, 24'd9116655, 24'd9004145, 24'd8769822, 24'd8460056, 24'd8136151, 24'd7862207, 24'd7692436, 24'd7660437, 24'd7772541, 24'd8006563, 24'd8316192, 24'd8640151, 24'd8914330, 24'd9084470, 24'd9116900, 24'd9005202, 24'd8771481, 
24'd8461990, 24'd8137977, 24'd7863563, 24'd7693055, 24'd7660195, 24'd7771486, 24'd8004905, 24'd8314258, 24'd8638324, 24'd8912972, 24'd9083849, 24'd9117139, 24'd9006254, 24'd8773138, 24'd8463924, 24'd8139805, 24'd7864923, 24'd7693678, 24'd7659958, 24'd7770436, 24'd8003249, 24'd8312324, 24'd8636496, 24'd8911610, 24'd9083224, 24'd9117374, 24'd9007302, 24'd8774792, 24'd8465857, 24'd8141634, 
24'd7866287, 24'd7694306, 24'd7659726, 24'd7769390, 24'd8001597, 24'd8310392, 24'd8634665, 24'd8910245, 24'd9082593, 24'd9117603, 24'd9008346, 24'd8776444, 24'd8467790, 24'd8143465, 24'd7867654, 24'd7694939, 24'd7659499, 24'd7768349, 24'd7999947, 24'd8308459, 24'd8632833, 24'd8908876, 24'd9081958, 24'd9117827, 24'd9009385, 24'd8778092, 24'd8469722, 24'd8145298, 24'd7869025, 24'd7695577, 
24'd7659278, 24'd7767312, 24'd7998299, 24'd8306528, 24'd8631000, 24'd8907503, 24'd9081317, 24'd9118046, 24'd9010420, 24'd8779739, 24'd8471653, 24'd8147133, 24'd7870400, 24'd7696220, 24'd7659061, 24'd7766279, 24'd7996655, 24'd8304597, 24'd8629164, 24'd8906126, 24'd9080672, 24'd9118260, 24'd9011451, 24'd8781382, 24'd8473584, 24'd8148969, 24'd7871778, 24'd7696867, 24'd7658850, 24'd7765251, 
24'd7995013, 24'd8302666, 24'd8627327, 24'd8904746, 24'd9080022, 24'd9118469, 24'd9012477, 24'd8783022, 24'd8475514, 24'd8150807, 24'd7873160, 24'd7697520, 24'd7658644, 24'd7764227, 24'd7993373, 24'd8300736, 24'd8625488, 24'd8903362, 24'd9079367, 24'd9118672, 24'd9013499, 24'd8784660, 24'd8477444, 24'd8152647, 24'd7874546, 24'd7698177, 24'd7658443, 24'd7763207, 24'd7991737, 24'd8298807, 
24'd8623648, 24'd8901975, 24'd9078708, 24'd9118871, 24'd9014516, 24'd8786295, 24'd8479372, 24'd8154488, 24'd7875935, 24'd7698839, 24'd7658247, 24'd7762192, 24'd7990104, 24'd8296878, 24'd8621806, 24'd8900584, 24'd9078043, 24'd9119064, 24'd9015529, 24'd8787927, 24'd8481301, 24'd8156331, 24'd7877328, 24'd7699506, 24'd7658056, 24'd7761181, 24'd7988473, 24'd8294950, 24'd8619962, 24'd8899190, 
24'd9077374, 24'd9119252, 24'd9016538, 24'd8789557, 24'd8483229, 24'd8158175, 24'd7878724, 24'd7700178, 24'd7657870, 24'd7760175, 24'd7986845, 24'd8293023, 24'd8618117, 24'd8897792, 24'd9076700, 24'd9119435, 24'd9017542, 24'd8791183, 24'd8485156, 24'd8160021, 24'd7880124, 24'd7700854, 24'd7657690, 24'd7759173, 24'd7985220, 24'd8291096, 24'd8616270, 24'd8896390, 24'd9076021, 24'd9119614, 
24'd9018542, 24'd8792807, 24'd8487082, 24'd8161869, 24'd7881527, 24'd7701536, 24'd7657514, 24'd7758175, 24'd7983597, 24'd8289170, 24'd8614422, 24'd8894985, 24'd9075337, 24'd9119786, 24'd9019537, 24'd8794428, 24'd8489008, 24'd8163718, 24'd7882934, 24'd7702222, 24'd7657344, 24'd7757182, 24'd7981978, 24'd8287245, 24'd8612571, 24'd8893576, 24'd9074648, 24'd9119954, 24'd9020528, 24'd8796046, 
24'd8490933, 24'd8165569, 24'd7884345, 24'd7702913, 24'd7657179, 24'd7756193, 24'd7980361, 24'd8285320, 24'd8610720, 24'd8892164, 24'd9073955, 24'd9120117, 24'd9021515, 24'd8797661, 24'd8492857, 24'd8167422, 24'd7885759, 24'd7703609, 24'd7657019, 24'd7755209, 24'd7978747, 24'd8283396, 24'd8608867, 24'd8890748, 24'd9073256, 24'd9120274, 24'd9022497, 24'd8799273, 24'd8494780, 24'd8169276, 
24'd7887176, 24'd7704309, 24'd7656864, 24'd7754229, 24'd7977136, 24'd8281473, 24'd8607012, 24'd8889328, 24'd9072553, 24'd9120427, 24'd9023474, 24'd8800883, 24'd8496703, 24'd8171131, 24'd7888598, 24'd7705015, 24'd7656714, 24'd7753253, 24'd7975528, 24'd8279551, 24'd8605155, 24'd8887906, 24'd9071846, 24'd9120574, 24'd9024448, 24'd8802490, 24'd8498625, 24'd8172988, 24'd7890022, 24'd7705725, 
24'd7656569, 24'd7752283, 24'd7973923, 24'd8277629, 24'd8603298, 24'd8886479, 24'd9071133, 24'd9120716, 24'd9025416, 24'd8804093, 24'd8500546, 24'd8174847, 24'd7891450, 24'd7706440, 24'd7656430, 24'd7751316, 24'd7972321, 24'd8275708, 24'd8601438, 24'd8885049, 24'd9070416, 24'd9120853, 24'd9026381, 24'd8805694, 24'd8502467, 24'd8176707, 24'd7892882, 24'd7707160, 24'd7656295, 24'd7750354, 
24'd7970722, 24'd8273788, 24'd8599577, 24'd8883616, 24'd9069693, 24'd9120985, 24'd9027340, 24'd8807292, 24'd8504386, 24'd8178568, 24'd7894317, 24'd7707885, 24'd7656166, 24'd7749396, 24'd7969125, 24'd8271869, 24'd8597715, 24'd8882179, 24'd9068966, 24'd9121112, 24'd9028296, 24'd8808887, 24'd8506305, 24'd8180432, 24'd7895755, 24'd7708614, 24'd7656042, 24'd7748443, 24'd7967532, 24'd8269951, 
24'd8595851, 24'd8880739, 24'd9068235, 24'd9121233, 24'd9029247, 24'd8810479, 24'd8508223, 24'd8182296, 24'd7897197, 24'd7709348, 24'd7655923, 24'd7747495, 24'd7965941, 24'd8268033, 24'd8593986, 24'd8879295, 24'd9067498, 24'd9121350, 24'd9030193, 24'd8812068, 24'd8510140, 24'd8184162, 24'd7898643, 24'd7710087, 24'd7655809, 24'd7746551, 24'd7964354, 24'd8266116, 24'd8592120, 24'd8877848, 
24'd9066757, 24'd9121461, 24'd9031135, 24'd8813654, 24'd8512057, 24'd8186029, 24'd7900092, 24'd7710831, 24'd7655700, 24'd7745611, 24'd7962769, 24'd8264200, 24'd8590251, 24'd8876397, 24'd9066011, 24'd9121567, 24'd9032072, 24'd8815237, 24'd8513972, 24'd8187898, 24'd7901544, 24'd7711579, 24'd7655597, 24'd7744676, 24'd7961188, 24'd8262285, 24'd8588382, 24'd8874943, 24'd9065260, 24'd9121668, 
24'd9033005, 24'd8816817, 24'd8515887, 24'd8189768, 24'd7903000, 24'd7712332, 24'd7655498, 24'd7743745, 24'd7959609, 24'd8260371, 24'd8586511, 24'd8873486, 24'd9064504, 24'd9121764, 24'd9033933, 24'd8818394, 24'd8517800, 24'd8191640, 24'd7904459, 24'd7713090, 24'd7655405, 24'd7742819, 24'd7958034, 24'd8258458, 24'd8584639, 24'd8872025, 24'd9063744, 24'd9121855, 24'd9034857, 24'd8819968, 
24'd8519713, 24'd8193513, 24'd7905921, 24'd7713853, 24'd7655317, 24'd7741898, 24'd7956461, 24'd8256546, 24'd8582765, 24'd8870561, 24'd9062979, 24'd9121940, 24'd9035776, 24'd8821539, 24'd8521625, 24'd8195387, 24'd7907387, 24'd7714620, 24'd7655234, 24'd7740981, 24'd7954892, 24'd8254634, 24'd8580890, 24'd8869093, 24'd9062209, 24'd9122021, 24'd9036691, 24'd8823107, 24'd8523536, 24'd8197263, 
24'd7908857, 24'd7715392, 24'd7655156, 24'd7740068, 24'd7953325, 24'd8252724, 24'd8579014, 24'd8867622, 24'd9061435, 24'd9122096, 24'd9037601, 24'd8824672, 24'd8525446, 24'd8199140, 24'd7910329, 24'd7716169, 24'd7655083, 24'd7739160, 24'd7951762, 24'd8250814, 24'd8577136, 24'd8866148, 24'd9060656, 24'd9122166, 24'd9038507, 24'd8826234, 24'd8527355, 24'd8201018, 24'd7911805, 24'd7716951, 
24'd7655015, 24'd7738257, 24'd7950201, 24'd8248906, 24'd8575257, 24'd8864670, 24'd9059872, 24'd9122231, 24'd9039408, 24'd8827793, 24'd8529263, 24'd8202898, 24'd7913285, 24'd7717737, 24'd7654953, 24'd7737358, 24'd7948644, 24'd8246998, 24'd8573377, 24'd8863189, 24'd9059083, 24'd9122291, 24'd9040305, 24'd8829348, 24'd8531170, 24'd8204779, 24'd7914767, 24'd7718528, 24'd7654896, 24'd7736464, 
24'd7947090, 24'd8245092, 24'd8571495, 24'd8861705, 24'd9058290, 24'd9122346, 24'd9041197, 24'd8830901, 24'd8533076, 24'd8206661, 24'd7916253, 24'd7719323, 24'd7654843, 24'd7735574, 24'd7945539, 24'd8243186, 24'd8569612, 24'd8860217, 24'd9057492, 24'd9122396, 24'd9042084, 24'd8832450, 24'd8534981, 24'd8208545, 24'd7917743, 24'd7720124, 24'd7654796, 24'd7734689, 24'd7943991, 24'd8241282, 
24'd8567728, 24'd8858726, 24'd9056689, 24'd9122440, 24'd9042967, 24'd8833997, 24'd8536885, 24'd8210430, 24'd7919235, 24'd7720929, 24'd7654755, 24'd7733809, 24'd7942446, 24'd8239378, 24'd8565842, 24'd8857232, 24'd9055882, 24'd9122480, 24'd9043845, 24'd8835540, 24'd8538788, 24'd8212316, 24'd7920731, 24'd7721738, 24'd7654718, 24'd7732933, 24'd7940904, 24'd8237476, 24'd8563956, 24'd8855735, 
24'd9055070, 24'd9122514, 24'd9044719, 24'd8837080, 24'd8540690, 24'd8214203, 24'd7922230, 24'd7722553, 24'd7654686, 24'd7732061, 24'd7939366, 24'd8235574, 24'd8562068, 24'd8854234, 24'd9054253, 24'd9122543, 24'd9045588, 24'd8838617, 24'd8542591, 24'd8216092, 24'd7923733, 24'd7723372, 24'd7654660, 24'd7731195, 24'd7937830, 24'd8233674, 24'd8560179, 24'd8852730, 24'd9053432, 24'd9122567, 
24'd9046452, 24'd8840151, 24'd8544491, 24'd8217981, 24'd7925238, 24'd7724195, 24'd7654638, 24'd7730332, 24'd7936298, 24'd8231775, 24'd8558288, 24'd8851222, 24'd9052606, 24'd9122585, 24'd9047312, 24'd8841682, 24'd8546390, 24'd8219872, 24'd7926747, 24'd7725024, 24'd7654622, 24'd7729475, 24'd7934769, 24'd8229877, 24'd8556397, 24'd8849712, 24'd9051775, 24'd9122599, 24'd9048167, 24'd8843210, 
24'd8548287, 24'd8221764, 24'd7928260, 24'd7725857, 24'd7654611, 24'd7728622, 24'd7933243, 24'd8227980, 24'd8554504, 24'd8848198, 24'd9050940, 24'd9122607, 24'd9049018, 24'd8844734, 24'd8550184, 24'd8223658, 24'd7929775, 24'd7726695, 24'd7654605, 24'd7727774, 24'd7931720, 24'd8226084, 24'd8552610, 24'd8846681, 24'd9050100, 24'd9122611, 24'd9049864, 24'd8846255, 24'd8552079, 24'd8225552, 
24'd7931294, 24'd7727537, 24'd7654605, 24'd7726930, 24'd7930201, 24'd8224189, 24'd8550715, 24'd8845161, 24'd9049255, 24'd9122609, 24'd9050705, 24'd8847773, 24'd8553973, 24'd8227448, 24'd7932816, 24'd7728384, 24'd7654609, 24'd7726091, 24'd7928684, 24'd8222295, 24'd8548819, 24'd8843637, 24'd9048406, 24'd9122602, 24'd9051541, 24'd8849288, 24'd8555866, 24'd8229344, 24'd7934341, 24'd7729235, 
24'd7654619, 24'd7725257, 24'd7927171, 24'd8220403, 24'd8546922, 24'd8842111, 24'd9047552, 24'd9122590, 24'd9052373, 24'd8850799, 24'd8557758, 24'd8231242, 24'd7935869, 24'd7730092, 24'd7654633, 24'd7724427, 24'd7925661, 24'd8218512, 24'd8545023, 24'd8840581, 24'd9046694, 24'd9122572, 24'd9053201, 24'd8852307, 24'd8559649, 24'd8233141, 24'd7937400, 24'd7730952, 24'd7654653, 24'd7723602, 
24'd7924155, 24'd8216621, 24'd8543124, 24'd8839048, 24'd9045831, 24'd9122550, 24'd9054023, 24'd8853812, 24'd8561538, 24'd8235041, 24'd7938935, 24'd7731818, 24'd7654678, 24'd7722782, 24'd7922651, 24'd8214733, 24'd8541223, 24'd8837512, 24'd9044963, 24'd9122522, 24'd9054841, 24'd8855314, 24'd8563426, 24'd8236942, 24'd7940472, 24'd7732688, 24'd7654708, 24'd7721966, 24'd7921151, 24'd8212845, 
24'd8539322, 24'd8835972, 24'd9044090, 24'd9122490, 24'd9055655, 24'd8856813, 24'd8565313, 24'd8238844, 24'd7942013, 24'd7733562, 24'd7654744, 24'd7721155, 24'd7919654, 24'd8210959, 24'd8537419, 24'd8834430, 24'd9043214, 24'd9122452, 24'd9056463, 24'd8858308, 24'd8567199, 24'd8240748, 24'd7943557, 24'd7734442, 24'd7654784, 24'd7720349, 24'd7918161, 24'd8209073, 24'd8535515, 24'd8832884, 
24'd9042332, 24'd9122409, 24'd9057267, 24'd8859800, 24'd8569084, 24'd8242652, 24'd7945104, 24'd7735325, 24'd7654830, 24'd7719547, 24'd7916671, 24'd8207189, 24'd8533611, 24'd8831336, 24'd9041446, 24'd9122361, 24'd9058067, 24'd8861288, 24'd8570967, 24'd8244557, 24'd7946655, 24'd7736214, 24'd7654880, 24'd7718750, 24'd7915184, 24'd8205307, 24'd8531705, 24'd8829784, 24'd9040555, 24'd9122307, 
24'd9058861, 24'd8862773, 24'd8572849, 24'd8246463, 24'd7948208, 24'd7737107, 24'd7654936, 24'd7717958, 24'd7913700, 24'd8203425, 24'd8529798, 24'd8828229, 24'd9039660, 24'd9122249, 24'd9059651, 24'd8864255, 24'd8574730, 24'd8248371, 24'd7949764, 24'd7738004, 24'd7654997, 24'd7717171, 24'd7912220, 24'd8201545, 24'd8527890, 24'd8826671, 24'd9038760, 24'd9122185, 24'd9060436, 24'd8865734, 
24'd8576609, 24'd8250279, 24'd7951324, 24'd7738906, 24'd7655064, 24'd7716388, 24'd7910743, 24'd8199667, 24'd8525981, 24'd8825110, 24'd9037856, 24'd9122116, 24'd9061217, 24'd8867209, 24'd8578487, 24'd8252188, 24'd7952886, 24'd7739813, 24'd7655135, 24'd7715610, 24'd7909269, 24'd8197789, 24'd8524072, 24'd8823546, 24'd9036947, 24'd9122043, 24'd9061993, 24'd8868681, 24'd8580364, 24'd8254098, 
24'd7954452, 24'd7740724, 24'd7655211, 24'd7714836, 24'd7907799, 24'd8195913, 24'd8522161, 24'd8821979, 24'd9036033, 24'd9121964, 24'd9062764, 24'd8870150, 24'd8582239, 24'd8256010, 24'd7956021, 24'd7741640, 24'd7655293, 24'd7714067, 24'd7906332, 24'd8194038, 24'd8520249, 24'd8820409, 24'd9035115, 24'd9121879, 24'd9063530, 24'd8871615, 24'd8584113, 24'd8257922, 24'd7957592, 24'd7742560, 
24'd7655380, 24'd7713303, 24'd7904869, 24'd8192165, 24'd8518337, 24'd8818836, 24'd9034193, 24'd9121790, 24'd9064292, 24'd8873077, 24'd8585986, 24'd8259835, 24'd7959167, 24'd7743485, 24'd7655472, 24'd7712544, 24'd7903409, 24'd8190293, 24'd8516424, 24'd8817259, 24'd9033266, 24'd9121696, 24'd9065049, 24'd8874535, 24'd8587857, 24'd8261749, 24'd7960745, 24'd7744414, 24'd7655569, 24'd7711790, 
24'd7901952, 24'd8188422, 24'd8514509, 24'd8815680, 24'd9032334, 24'd9121596, 24'd9065801, 24'd8875990, 24'd8589727, 24'd8263663, 24'd7962326, 24'd7745348, 24'd7655671, 24'd7711040, 24'd7900499, 24'd8186553, 24'd8512594, 24'd8814098, 24'd9031398, 24'd9121491, 24'd9066548, 24'd8877442, 24'd8591596, 24'd8265579, 24'd7963909, 24'd7746287, 24'd7655778, 24'd7710295, 24'd7899049, 24'd8184686, 
24'd8510678, 24'd8812513, 24'd9030458, 24'd9121381, 24'd9067291, 24'd8878890, 24'd8593463, 24'd8267495, 24'd7965496, 24'd7747229, 24'd7655890, 24'd7709555, 24'd7897603, 24'd8182819, 24'd8508761, 24'd8810925, 24'd9029512, 24'd9121266, 24'd9068029, 24'd8880334, 24'd8595328, 24'd8269413, 24'd7967086, 24'd7748177, 24'd7656008, 24'd7708819, 24'd7896160, 24'd8180954, 24'd8506843, 24'd8809333, 
24'd9028563, 24'd9121146, 24'd9068762, 24'd8881776, 24'd8597193, 24'd8271331, 24'd7968678, 24'd7749129, 24'd7656131, 24'd7708089, 24'd7894720, 24'd8179091, 24'd8504925, 24'd8807739, 24'd9027609, 24'd9121021, 24'd9069490, 24'd8883213, 24'd8599055, 24'd8273250, 24'd7970274, 24'd7750085, 24'd7656259, 24'd7707363, 24'd7893284, 24'd8177229, 24'd8503005, 24'd8806142, 24'd9026650, 24'd9120891, 
24'd9070213, 24'd8884648, 24'd8600917, 24'd8275170, 24'd7971872, 24'd7751046, 24'd7656392, 24'd7706642, 24'd7891851, 24'd8175368, 24'd8501085, 24'd8804542, 24'd9025687, 24'd9120755, 24'd9070932, 24'd8886079, 24'd8602776, 24'd8277090, 24'd7973474, 24'd7752011, 24'd7656530, 24'd7705925, 24'd7890422, 24'd8173509, 24'd8499164, 24'd8802940, 24'd9024720, 24'd9120614, 24'd9071646, 24'd8887506, 
24'd8604635, 24'd8279012, 24'd7975078, 24'd7752981, 24'd7656673, 24'd7705214, 24'd7888997, 24'd8171652, 24'd8497242, 24'd8801334, 24'd9023748, 24'd9120469, 24'd9072355, 24'd8888930, 24'd8606491, 24'd8280934, 24'd7976685, 24'd7753955, 24'd7656821, 24'd7704507, 24'd7887575, 24'd8169796, 24'd8495320, 24'd8799725, 24'd9022771, 24'd9120318, 24'd9073060, 24'd8890350, 24'd8608347, 24'd8282857, 
24'd7978295, 24'd7754934, 24'd7656975, 24'd7703805, 24'd7886156, 24'd8167941, 24'd8493396, 24'd8798114, 24'd9021790, 24'd9120162, 24'd9073759, 24'd8891767, 24'd8610200, 24'd8284781, 24'd7979908, 24'd7755917, 24'd7657133, 24'd7703108, 24'd7884741, 24'd8166089, 24'd8491472, 24'd8796499, 24'd9020805, 24'd9120000, 24'd9074454, 24'd8893180, 24'd8612052, 24'd8286705, 24'd7981524, 24'd7756904, 
24'd7657297, 24'd7702415, 24'd7883329, 24'd8164237, 24'd8489547, 24'd8794882, 24'd9019815, 24'd9119834, 24'd9075144, 24'd8894590, 24'd8613903, 24'd8288630, 24'd7983143, 24'd7757896, 24'd7657466, 24'd7701728, 24'd7881921, 24'd8162387, 24'd8487622, 24'd8793262, 24'd9018821, 24'd9119663, 24'd9075829, 24'd8895996, 24'd8615752, 24'd8290556, 24'd7984764, 24'd7758892, 24'd7657640, 24'd7701045, 
24'd7880517, 24'd8160539, 24'd8485696, 24'd8791639, 24'd9017823, 24'd9119486, 24'd9076510, 24'd8897399, 24'd8617599, 24'd8292482, 24'd7986389, 24'd7759893, 24'd7657819, 24'd7700367, 24'd7879116, 24'd8158693, 24'd8483769, 24'd8790013, 24'd9016820, 24'd9119304, 24'd9077185, 24'd8898798, 24'd8619445, 24'd8294410, 24'd7988016, 24'd7760898, 24'd7658004, 24'd7699694, 24'd7877719, 24'd8156848, 
24'd8481842, 24'd8788384, 24'd9015812, 24'd9119117, 24'd9077856, 24'd8900194, 24'd8621289, 24'd8296337, 24'd7989646, 24'd7761908, 24'd7658193, 24'd7699026, 24'd7876325, 24'd8155004, 24'd8479913, 24'd8786753, 24'd9014800, 24'd9118925, 24'd9078522, 24'd8901585, 24'd8623132, 24'd8298266, 24'd7991279, 24'd7762922, 24'd7658387, 24'd7698362, 24'd7874935, 24'd8153163, 24'd8477985, 24'd8785119, 
24'd9013784, 24'd9118728, 24'd9079183, 24'd8902974, 24'd8624973, 24'd8300195, 24'd7992914, 24'd7763940, 24'd7658587, 24'd7697703, 24'd7873548, 24'd8151323, 24'd8476055, 24'd8783482, 24'd9012764, 24'd9118526, 24'd9079839, 24'd8904358, 24'd8626812, 24'd8302125, 24'd7994553, 24'd7764963, 24'd7658792, 24'd7697050, 24'd7872166, 24'd8149484, 24'd8474125, 24'd8781842, 24'd9011739, 24'd9118319, 
24'd9080490, 24'd8905740, 24'd8628649, 24'd8304055, 24'd7996194, 24'd7765990, 24'd7659002, 24'd7696401, 24'd7870786, 24'd8147648, 24'd8472194, 24'd8780200, 24'd9010709, 24'd9118106, 24'd9081137, 24'd8907117, 24'd8630485, 24'd8305986, 24'd7997838, 24'd7767022, 24'd7659217, 24'd7695757, 24'd7869411, 24'd8145813, 24'd8470263, 24'd8778554, 24'd9009676, 24'd9117889, 24'd9081779, 24'd8908491, 
24'd8632319, 24'd8307918, 24'd7999484, 24'd7768058, 24'd7659437, 24'd7695117, 24'd7868039, 24'd8143979, 24'd8468331, 24'd8776906, 24'd9008638, 24'd9117666, 24'd9082415, 24'd8909861, 24'd8634152, 24'd8309850, 24'd8001134, 24'd7769098, 24'd7659662, 24'd7694483, 24'd7866670, 24'd8142148, 24'd8466399, 24'd8775256, 24'd9007595, 24'd9117438, 24'd9083047, 24'd8911228, 24'd8635983, 24'd8311782, 
24'd8002786, 24'd7770142, 24'd7659892, 24'd7693854, 24'd7865305, 24'd8140318, 24'd8464466, 24'd8773602, 24'd9006549, 24'd9117206, 24'd9083674, 24'd8912591, 24'd8637812, 24'd8313715, 24'd8004440, 24'd7771191, 24'd7660128, 24'd7693229, 24'd7863944, 24'd8138490, 24'd8462533, 24'd8771946, 24'd9005498, 24'd9116968, 24'd9084296, 24'd8913950, 24'd8639639, 24'd8315649, 24'd8006098, 24'd7772245, 
24'd7660368, 24'd7692609, 24'd7862587, 24'd8136663, 24'd8460599, 24'd8770287, 24'd9004442, 24'd9116724, 24'd9084914, 24'd8915305, 24'd8641464, 24'd8317583, 24'd8007758, 24'd7773302, 24'd7660614, 24'd7691994, 24'd7861233, 24'd8134839, 24'd8458664, 24'd8768626, 24'd9003383, 24'd9116476, 24'd9085526, 24'd8916657, 24'd8643288, 24'd8319518, 24'd8009421, 24'd7774364, 24'd7660865, 24'd7691384, 
24'd7859883, 24'd8133016, 24'd8456729, 24'd8766962, 24'd9002319, 24'd9116223, 24'd9086134, 24'd8918005, 24'd8645110, 24'd8321453, 24'd8011086, 24'd7775430, 24'd7661121, 24'd7690779, 24'd7858537, 24'd8131195, 24'd8454794, 24'd8765295, 24'd9001250, 24'd9115965, 24'd9086736, 24'd8919350, 24'd8646930, 24'd8323389, 24'd8012754, 24'd7776501, 24'd7661382, 24'd7690179, 24'd7857195, 24'd8129376, 
24'd8452858, 24'd8763626, 24'd9000178, 24'd9115701, 24'd9087334, 24'd8920690, 24'd8648748, 24'd8325325, 24'd8014425, 24'd7777575, 24'd7661648, 24'd7689584, 24'd7855856, 24'd8127558, 24'd8450922, 24'd8761953, 24'd8999101, 24'd9115432, 24'd9087927, 24'd8922027, 24'd8650565, 24'd8327262, 24'd8016099, 24'd7778654, 24'd7661919, 24'd7688994, 24'd7854521, 24'd8125743, 24'd8448985, 24'd8760279, 
24'd8998020, 24'd9115159, 24'd9088515, 24'd8923361, 24'd8652380, 24'd8329199, 24'd8017775, 24'd7779738, 24'd7662195, 24'd7688408, 24'd7853189, 24'd8123929, 24'd8447048, 24'd8758601, 24'd8996934, 24'd9114880, 24'd9089098, 24'd8924690, 24'd8654192, 24'd8331136, 24'd8019453, 24'd7780825, 24'd7662476, 24'd7687827, 24'd7851862, 24'd8122117, 24'd8445110, 24'd8756922, 24'd8995844, 24'd9114596, 
24'd9089676, 24'd8926016, 24'd8656003, 24'd8333074, 24'd8021134, 24'd7781917, 24'd7662763, 24'd7687252, 24'd7850538, 24'd8120307, 24'd8443172, 24'd8755239, 24'd8994750, 24'd9114307, 24'd9090249, 24'd8927338, 24'd8657812, 24'd8335012, 24'd8022818, 24'd7783013, 24'd7663054, 24'd7686681, 24'd7849218, 24'd8118499, 24'd8441234, 24'd8753554, 24'd8993652, 24'd9114013, 24'd9090817, 24'd8928656, 
24'd8659620, 24'd8336951, 24'd8024504, 24'd7784114, 24'd7663351, 24'd7686115, 24'd7847902, 24'd8116693, 24'd8439295, 24'd8751867, 24'd8992550, 24'd9113714, 24'd9091381, 24'd8929970, 24'd8661425, 24'd8338890, 24'd8026193, 24'd7785218, 24'd7663653, 24'd7685554, 24'd7846589, 24'd8114888, 24'd8437356, 24'd8750176, 24'd8991443, 24'd9113410, 24'd9091939, 24'd8931281, 24'd8663228, 24'd8340829, 
24'd8027885, 24'd7786327, 24'd7663959, 24'd7684998, 24'd7845280, 24'd8113086, 24'd8435416, 24'd8748484, 24'd8990332, 24'd9113100, 24'd9092493, 24'd8932588, 24'd8665030, 24'd8342768, 24'd8029579, 24'd7787440, 24'd7664271, 24'd7684447, 24'd7843975, 24'd8111285, 24'd8433477, 24'd8746788, 24'd8989217, 24'd9112786, 24'd9093041, 24'd8933891, 24'd8666829, 24'd8344708, 24'd8031275, 24'd7788557, 
24'd7664588, 24'd7683901, 24'd7842674, 24'd8109487, 24'd8431537, 24'd8745091, 24'd8988098, 24'd9112466, 24'd9093585, 24'd8935190, 24'd8668627, 24'd8346649, 24'd8032974, 24'd7789679, 24'd7664910, 24'd7683360, 24'd7841377, 24'd8107690, 24'd8429596, 24'd8743391, 24'd8986974, 24'd9112142, 24'd9094124, 24'd8936485, 24'd8670422, 24'd8348589, 24'd8034675, 24'd7790804, 24'd7665237, 24'd7682824, 
24'd7840084, 24'd8105896, 24'd8427655, 24'd8741688, 24'd8985846, 24'd9111812, 24'd9094657, 24'd8937776, 24'd8672216, 24'd8350530, 24'd8036379, 24'd7791934, 24'd7665569, 24'd7682293, 24'd7838794, 24'd8104103, 24'd8425714, 24'd8739983, 24'd8984714, 24'd9111478, 24'd9095186, 24'd8939064, 24'd8674008, 24'd8352471, 24'd8038086, 24'd7793068, 24'd7665907, 24'd7681766, 24'd7837509, 24'd8102312, 
24'd8423773, 24'd8738275, 24'd8983578, 24'd9111138, 24'd9095710, 24'd8940348, 24'd8675797, 24'd8354412, 24'd8039795, 24'd7794206, 24'd7666249, 24'd7681245, 24'd7836227, 24'd8100524, 24'd8421832, 24'd8736565, 24'd8982438, 24'd9110793, 24'd9096229, 24'd8941628, 24'd8677585, 24'd8356354, 24'd8041506, 24'd7795349, 24'd7666596, 24'd7680729, 24'd7834949, 24'd8098737, 24'd8419890, 24'd8734852, 
24'd8981294, 24'd9110443, 24'd9096743, 24'd8942904, 24'd8679371, 24'd8358296, 24'd8043220, 24'd7796495, 24'd7666949, 24'd7680217, 24'd7833675, 24'd8096952, 24'd8417948, 24'd8733137, 24'd8980145, 24'd9110088, 24'd9097252, 24'd8944176, 24'd8681154, 24'd8360238, 24'd8044936, 24'd7797646, 24'd7667306, 24'd7679711, 24'd7832404, 24'd8095170, 24'd8416006, 24'd8731420, 24'd8978992, 24'd9109728, 
24'd9097756, 24'd8945444, 24'd8682936, 24'd8362180, 24'd8046654, 24'd7798801, 24'd7667669, 24'd7679209, 24'd7831138, 24'd8093389, 24'd8414064, 24'd8729700, 24'd8977835, 24'd9109363, 24'd9098255, 24'd8946708, 24'd8684715, 24'd8364122, 24'd8048375, 24'd7799960, 24'd7668036, 24'd7678713, 24'd7829876, 24'd8091611, 24'd8412121, 24'd8727978, 24'd8976674, 24'd9108993, 24'd9098749, 24'd8947969, 
24'd8686492, 24'd8366065, 24'd8050099, 24'd7801123, 24'd7668409, 24'd7678221, 24'd7828617, 24'd8089835, 24'd8410179, 24'd8726254, 24'd8975509, 24'd9108618, 24'd9099238, 24'd8949225, 24'd8688268, 24'd8368008, 24'd8051825, 24'd7802290, 24'd7668787, 24'd7677735, 24'd7827363, 24'd8088060, 24'd8408236, 24'd8724527, 24'd8974340, 24'd9108238, 24'd9099722, 24'd8950478, 24'd8690041, 24'd8369951, 
24'd8053553, 24'd7803461, 24'd7669169, 24'd7677253, 24'd7826112, 24'd8086288, 24'd8406293, 24'd8722797, 24'd8973166, 24'd9107852, 24'd9100201, 24'd8951727, 24'd8691812, 24'd8371894, 24'd8055283, 24'd7804637, 24'd7669557, 24'd7676776, 24'd7824866, 24'd8084518, 24'd8404350, 24'd8721066, 24'd8971989, 24'd9107462, 24'd9100675, 24'd8952971, 24'd8693581, 24'd8373837, 24'd8057016, 24'd7805816, 
24'd7669950, 24'd7676305, 24'd7823623, 24'd8082750, 24'd8402407, 24'd8719332, 24'd8970807, 24'd9107067, 24'd9101144, 24'd8954212, 24'd8695348, 24'd8375780, 24'd8058751, 24'd7807000, 24'd7670348, 24'd7675838, 24'd7822384, 24'd8080985, 24'd8400463, 24'd8717596, 24'd8969622, 24'd9106666, 24'd9101608, 24'd8955449, 24'd8697112, 24'd8377723, 24'd8060488, 24'd7808188, 24'd7670751, 24'd7675377, 
24'd7821149, 24'd8079221, 24'd8398520, 24'd8715857, 24'd8968432, 24'd9106261, 24'd9102067, 24'd8956681, 24'd8698875, 24'd8379667, 24'd8062228, 24'd7809379, 24'd7671159, 24'd7674920, 24'd7819919, 24'd8077460, 24'd8396577, 24'd8714116, 24'd8967238, 24'd9105850, 24'd9102521, 24'd8957910, 24'd8700635, 24'd8381610, 24'd8063970, 24'd7810575, 24'd7671572, 24'd7674468, 24'd7818692, 24'd8075701, 
24'd8394633, 24'd8712373, 24'd8966040, 24'd9105435, 24'd9102971, 24'd8959135, 24'd8702393, 24'd8383554, 24'd8065714, 24'd7811775, 24'd7671990, 24'd7674022, 24'd7817469, 24'd8073944, 24'd8392689, 24'd8710628, 24'd8964839, 24'd9105014, 24'd9103415, 24'd8960356, 24'd8704149, 24'd8385497, 24'd8067461, 24'd7812979, 24'd7672413, 24'd7673580, 24'd7816250, 24'd8072189, 24'd8390746, 24'd8708880, 
24'd8963633, 24'd9104589, 24'd9103854, 24'd8961573, 24'd8705903, 24'd8387441, 24'd8069210, 24'd7814187, 24'd7672841, 24'd7673144, 24'd7815035, 24'd8070436, 24'd8388802, 24'd8707130, 24'd8962423, 24'd9104158, 24'd9104288, 24'd8962785, 24'd8707654, 24'd8389384, 24'd8070961, 24'd7815399, 24'd7673274, 24'd7672712, 24'd7813825, 24'd8068686, 24'd8386859, 24'd8705378, 24'd8961209, 24'd9103723, 
24'd9104717, 24'd8963994, 24'd8709404, 24'd8391328, 24'd8072714, 24'd7816615, 24'd7673712, 24'd7672285, 24'd7812618, 24'd8066938, 24'd8384915, 24'd8703623, 24'd8959991, 24'd9103282, 24'd9105141, 24'd8965199, 24'd8711151, 24'd8393272, 24'd8074470, 24'd7817835, 24'd7674155, 24'd7671864, 24'd7811415, 24'd8065192, 24'd8382972, 24'd8701867, 24'd8958769, 24'd9102837, 24'd9105560, 24'd8966400, 
24'd8712895, 24'd8395215, 24'd8076227, 24'd7819059, 24'd7674603, 24'd7671447, 24'd7810217, 24'd8063448, 24'd8381028, 24'd8700108, 24'd8957543, 24'd9102386, 24'd9105974, 24'd8967596, 24'd8714638, 24'd8397159, 24'd8077987, 24'd7820287, 24'd7675056, 24'd7671036, 24'd7809022, 24'd8061707, 24'd8379085, 24'd8698347, 24'd8956313, 24'd9101930, 24'd9106383, 24'd8968789, 24'd8716378, 24'd8399102, 
24'd8079749, 24'd7821519, 24'd7675514, 24'd7670630, 24'd7807831, 24'd8059968, 24'd8377141, 24'd8696584, 24'd8955079, 24'd9101470, 24'd9106787, 24'd8969977, 24'd8718116, 24'd8401045, 24'd8081513, 24'd7822755, 24'd7675977, 24'd7670228, 24'd7806645, 24'd8058231, 24'd8375198, 24'd8694819, 24'd8953841, 24'd9101004, 24'd9107186, 24'd8971162, 24'd8719851, 24'd8402989, 24'd8083280, 24'd7823995, 
24'd7676445, 24'd7669832, 24'd7805463, 24'd8056497, 24'd8373255, 24'd8693051, 24'd8952599, 24'd9100534, 24'd9107579, 24'd8972342, 24'd8721585, 24'd8404932, 24'd8085048, 24'd7825239, 24'd7676919, 24'd7669441, 24'd7804284, 24'd8054765, 24'd8371312, 24'd8691282, 24'd8951353, 24'd9100058, 24'd9107968, 24'd8973518, 24'd8723316, 24'd8406875, 24'd8086819, 24'd7826486, 24'd7677397, 24'd7669054, 
24'd7803110, 24'd8053035, 24'd8369369, 24'd8689510, 24'd8950103, 24'd9099577, 24'd9108352, 24'd8974690, 24'd8725044, 24'd8408818, 24'd8088592, 24'd7827738, 24'd7677880, 24'd7668673, 24'd7801940, 24'd8051307, 24'd8367426, 24'd8687736, 24'd8948849, 24'd9099092, 24'd9108731, 24'd8975858, 24'd8726770, 24'd8410760, 24'd8090366, 24'd7828994, 24'd7678368, 24'd7668297, 24'd7800774, 24'd8049582, 
24'd8365483, 24'd8685960, 24'd8947592, 24'd9098601, 24'd9109104, 24'd8977022, 24'd8728494, 24'd8412703, 24'd8092143, 24'd7830254, 24'd7678861, 24'd7667926, 24'd7799612, 24'd8047860, 24'd8363541, 24'd8684182, 24'd8946330, 24'd9098106, 24'd9109473, 24'd8978182, 24'd8730216, 24'd8414645, 24'd8093922, 24'd7831517, 24'd7679359, 24'd7667560, 24'd7798454, 24'd8046140, 24'd8361598, 24'd8682402, 
24'd8945065, 24'd9097605, 24'd9109837, 24'd8979338, 24'd8731935, 24'd8416588, 24'd8095704, 24'd7832785, 24'd7679862, 24'd7667199, 24'd7797301, 24'd8044422, 24'd8359656, 24'd8680620, 24'd8943795, 24'd9097100, 24'd9110195, 24'd8980489, 24'd8733651, 24'd8418530, 24'd8097487, 24'd7834056, 24'd7680370, 24'd7666843, 24'd7796151, 24'd8042706, 24'd8357714, 24'd8678836, 24'd8942522, 24'd9096589, 
24'd9110548, 24'd8981637, 24'd8735366, 24'd8420472, 24'd8099272, 24'd7835331, 24'd7680883, 24'd7666492, 24'd7795006, 24'd8040993, 24'd8355772, 24'd8677050, 24'd8941245, 24'd9096074, 24'd9110897, 24'd8982780, 24'd8737077, 24'd8422413, 24'd8101059, 24'd7836610, 24'd7681401, 24'd7666146, 24'd7793865, 24'd8039283, 24'd8353831, 24'd8675262, 24'd8939964, 24'd9095554, 24'd9111240, 24'd8983919, 
24'd8738787, 24'd8424355, 24'd8102848, 24'd7837893, 24'd7681923, 24'd7665805, 24'd7792728, 24'd8037574, 24'd8351890, 24'd8673471, 24'd8938679, 24'd9095028, 24'd9111578, 24'd8985054, 24'd8740494, 24'd8426296, 24'd8104640, 24'd7839180, 24'd7682451, 24'd7665469, 24'd7791595, 24'd8035869, 24'd8349949, 24'd8671679, 24'd8937390, 24'd9094498, 24'd9111912, 24'd8986185, 24'd8742198, 24'd8428237, 
24'd8106433, 24'd7840471, 24'd7682984, 24'd7665139, 24'd7790467, 24'd8034166, 24'd8348008, 24'd8669885, 24'd8936097, 24'd9093963, 24'd9112240, 24'd8987311, 24'd8743900, 24'd8430177, 24'd8108228, 24'd7841765, 24'd7683522, 24'd7664813, 24'd7789342, 24'd8032465, 24'd8346067, 24'd8668089, 24'd8934801, 24'd9093423, 24'd9112563, 24'd8988433, 24'd8745600, 24'd8432118, 24'd8110025, 24'd7843064, 
24'd7684064, 24'd7664493, 24'd7788222, 24'd8030767, 24'd8344127, 24'd8666290, 24'd8933501, 24'd9092878, 24'd9112881, 24'd8989551, 24'd8747296, 24'd8434058, 24'd8111824, 24'd7844366, 24'd7684612, 24'd7664177, 24'd7787106, 24'd8029071, 24'd8342187, 24'd8664490, 24'd8932197, 24'd9092328, 24'd9113194, 24'd8990665, 24'd8748991, 24'd8435997, 24'd8113625, 24'd7845672, 24'd7685164, 24'd7663867, 
24'd7785994, 24'd8027378, 24'd8340248, 24'd8662688, 24'd8930889, 24'd9091773, 24'd9113501, 24'd8991775, 24'd8750683, 24'd8437937, 24'd8115428, 24'd7846982, 24'd7685722, 24'd7663562, 24'd7784887, 24'd8025687, 24'd8338309, 24'd8660884, 24'd8929577, 24'd9091213, 24'd9113804, 24'd8992880, 24'd8752372, 24'd8439876, 24'd8117233, 24'd7848295, 24'd7686284, 24'd7663262, 24'd7783784, 24'd8023999, 
24'd8336370, 24'd8659079, 24'd8928261, 24'd9090648, 24'd9114102, 24'd8993982, 24'd8754059, 24'd8441814, 24'd8119040, 24'd7849613, 24'd7686851, 24'd7662966, 24'd7782684, 24'd8022314, 24'd8334431, 24'd8657271, 24'd8926942, 24'd9090078, 24'd9114394, 24'd8995079, 24'd8755743, 24'd8443753, 24'd8120849, 24'd7850934, 24'd7687424, 24'd7662676, 24'd7781590, 24'd8020631, 24'd8332493, 24'd8655461, 
24'd8925619, 24'd9089503, 24'd9114682, 24'd8996171, 24'd8757425, 24'd8445691, 24'd8122659, 24'd7852259, 24'd7688001, 24'd7662392, 24'd7780499, 24'd8018950, 24'd8330556, 24'd8653650, 24'd8924292, 24'd9088924, 24'd9114964, 24'd8997260, 24'd8759104, 24'd8447628, 24'd8124472, 24'd7853588, 24'd7688583, 24'd7662112, 24'd7779413, 24'd8017272, 24'd8328618, 24'd8651836, 24'd8922962, 24'd9088339, 
24'd9115241, 24'd8998344, 24'd8760781, 24'd8449565, 24'd8126286, 24'd7854920, 24'd7689170, 24'd7661837, 24'd7778331, 24'd8015597, 24'd8326682, 24'd8650021, 24'd8921627, 24'd9087750, 24'd9115513, 24'd8999424, 24'd8762455, 24'd8451502, 24'd8128102, 24'd7856256, 24'd7689762, 24'd7661567, 24'd7777253, 24'd8013925, 24'd8324745, 24'd8648204, 24'd8920289, 24'd9087156, 24'd9115781, 24'd9000499, 
24'd8764126, 24'd8453438, 24'd8129920, 24'd7857596, 24'd7690358, 24'd7661303, 24'd7776180, 24'd8012255, 24'd8322809, 24'd8646385, 24'd8918947, 24'd9086556, 24'd9116043, 24'd9001571, 24'd8765794, 24'd8455374, 24'd8131740, 24'd7858940, 24'd7690960, 24'd7661043, 24'd7775110, 24'd8010587, 24'd8320874, 24'd8644564, 24'd8917602, 24'd9085952, 24'd9116299, 24'd9002638, 24'd8767460, 24'd8457309, 
24'd8133562, 24'd7860287, 24'd7691567, 24'd7660789, 24'd7774045, 24'd8008923, 24'd8318939, 24'd8642742, 24'd8916253, 24'd9085343, 24'd9116551, 24'd9003700, 24'd8769124, 24'd8459244, 24'd8135385, 24'd7861638, 24'd7692178, 24'd7660540, 24'd7772985, 24'd8007261, 24'd8317004, 24'd8640918, 24'd8914900, 24'd9084729, 24'd9116798, 24'd9004759, 24'd8770784, 24'd8461178, 24'd8137210, 24'd7862993, 
24'd7692794, 24'd7660296, 24'd7771929, 24'd8005601, 24'd8315070, 24'd8639092, 24'd8913543, 24'd9084111, 24'd9117039, 24'd9005813, 24'd8772442, 24'd8463112, 24'd8139037, 24'd7864352, 24'd7693416, 24'd7660057, 24'd7770877, 24'd8003945, 24'd8313136, 24'd8637264, 24'd8912183, 24'd9083487, 24'd9117276, 24'd9006863, 24'd8774098, 24'd8465045, 24'd8140866, 24'd7865714, 24'd7694042, 24'd7659823, 
24'd7769829, 24'd8002291, 24'd8311203, 24'd8635434, 24'd8910819, 24'd9082858, 24'd9117507, 24'd9007908, 24'd8775750, 24'd8466978, 24'd8142696, 24'd7867080, 24'd7694673, 24'd7659594, 24'd7768786, 24'd8000639, 24'd8309271, 24'd8633603, 24'd8909451, 24'd9082225, 24'd9117733, 24'd9008949, 24'd8777400, 24'd8468910, 24'd8144528, 24'd7868449, 24'd7695308, 24'd7659370, 24'd7767747, 24'd7998991, 
24'd8307339, 24'd8631770, 24'd8908080, 24'd9081587, 24'd9117955, 24'd9009986, 24'd8779047, 24'd8470842, 24'd8146362, 24'd7869822, 24'd7695949, 24'd7659152, 24'd7766712, 24'd7997345, 24'd8305408, 24'd8629935, 24'd8906705, 24'd9080944, 24'd9118171, 24'd9011018, 24'd8780692, 24'd8472773, 24'd8148197, 24'd7871199, 24'd7696595, 24'd7658938, 24'd7765682, 24'd7995702, 24'd8303477, 24'd8628099, 
24'd8905326, 24'd9080296, 24'd9118381, 24'd9012046, 24'd8782334, 24'd8474703, 24'd8150035, 24'd7872579, 24'd7697245, 24'd7658730, 24'd7764656, 24'd7994062, 24'd8301547, 24'd8626261, 24'd8903944, 24'd9079643, 24'd9118587, 24'd9013070, 24'd8783972, 24'd8476633, 24'd8151874, 24'd7873963, 24'd7697900, 24'd7658527, 24'd7763635, 24'd7992424, 24'd8299617, 24'd8624421, 24'd8902558, 24'd9078985, 
24'd9118788, 24'd9014089, 24'd8785609, 24'd8478562, 24'd8153714, 24'd7875351, 24'd7698560, 24'd7658329, 24'd7762618, 24'd7990789, 24'd8297688, 24'd8622580, 24'd8901169, 24'd9078323, 24'd9118983, 24'd9015104, 24'd8787242, 24'd8480491, 24'd8155556, 24'd7876742, 24'd7699225, 24'd7658136, 24'd7761605, 24'd7989157, 24'd8295760, 24'd8620737, 24'd8899776, 24'd9077656, 24'd9119174, 24'd9016114, 
24'd8788873, 24'd8482419, 24'd8157400, 24'd7878137, 24'd7699895, 24'd7657948, 24'd7760597, 24'd7987528, 24'd8293832, 24'd8618892, 24'd8898379, 24'd9076983, 24'd9119359, 24'd9017121, 24'd8790500, 24'd8484346, 24'd8159246, 24'd7879535, 24'd7700569, 24'd7657765, 24'd7759593, 24'd7985902, 24'd8291905, 24'd8617046, 24'd8896979, 24'd9076306, 24'd9119539, 24'd9018122, 24'd8792125, 24'd8486273, 
24'd8161093, 24'd7880937, 24'd7701249, 24'd7657587, 24'd7758594, 24'd7984278, 24'd8289979, 24'd8615198, 24'd8895575, 24'd9075625, 24'd9119714, 24'd9019119, 24'd8793747, 24'd8488199, 24'd8162941, 24'd7882343, 24'd7701933, 24'd7657415, 24'd7757599, 24'd7982658, 24'd8288054, 24'd8613349, 24'd8894168, 24'd9074938, 24'd9119884, 24'd9020112, 24'd8795367, 24'd8490124, 24'd8164792, 24'd7883752, 
24'd7702622, 24'd7657248, 24'd7756608, 24'd7981040, 24'd8286129, 24'd8611498, 24'd8892757, 24'd9074247, 24'd9120049, 24'd9021101, 24'd8796983, 24'd8492049, 24'd8166643, 24'd7885164, 24'd7703316, 24'd7657085, 24'd7755622, 24'd7979425, 24'd8284204, 24'd8609645, 24'd8891343, 24'd9073550, 24'd9120209, 24'd9022085, 24'd8798597, 24'd8493972, 24'd8168497, 24'd7886580, 24'd7704015, 24'd7656928, 
24'd7754640, 24'd7977813, 24'd8282281, 24'd8607791, 24'd8889925, 24'd9072849, 24'd9120363, 24'd9023064, 24'd8800207, 24'd8495895, 24'd8170352, 24'd7888000, 24'd7704718, 24'd7656776, 24'd7753663, 24'd7976203, 24'd8280358, 24'd8605935, 24'd8888504, 24'd9072144, 24'd9120513, 24'd9024039, 24'd8801815, 24'd8497818, 24'd8172208, 24'd7889423, 24'd7705426, 24'd7656629, 24'd7752690, 24'd7974597, 
24'd8278436, 24'd8604078, 24'd8887079, 24'd9071433, 24'd9120657, 24'd9025010, 24'd8803420, 24'd8499739, 24'd8174066, 24'd7890850, 24'd7706139, 24'd7656488, 24'd7751721, 24'd7972994, 24'd8276515, 24'd8602220, 24'd8885650, 24'd9070717, 24'd9120796, 24'd9025976, 24'd8805022, 24'd8501660, 24'd8175925, 24'd7892280, 24'd7706857, 24'd7656351, 24'd7750757, 24'd7971393, 24'd8274595, 24'd8600359, 
24'd8884219, 24'd9069997, 24'd9120930, 24'd9026938, 24'd8806621, 24'd8503580, 24'd8177786, 24'd7893714, 24'd7707580, 24'd7656220, 24'd7749798, 24'd7969796, 24'd8272675, 24'd8598498, 24'd8882783, 24'd9069272, 24'd9121059, 24'd9027895, 24'd8808217, 24'd8505499, 24'd8179649, 24'd7895151, 24'd7708307, 24'd7656093, 24'd7748843, 24'd7968201, 24'd8270756, 24'd8596634, 24'd8881344, 24'd9068543, 
24'd9121183, 24'd9028848, 24'd8809810, 24'd8507418, 24'd8181513, 24'd7896591, 24'd7709039, 24'd7655972, 24'd7747893, 24'd7966609, 24'd8268838, 24'd8594770, 24'd8879902, 24'd9067808, 24'd9121301, 24'd9029796, 24'd8811401, 24'd8509335, 24'd8183378, 24'd7898035, 24'd7709776, 24'd7655856, 24'd7746947, 24'd7965020, 24'd8266921, 24'd8592904, 24'd8878456, 24'd9067069, 24'd9121415, 24'd9030740, 
24'd8812988, 24'd8511252, 24'd8185245, 24'd7899483, 24'd7710518, 24'd7655745, 24'd7746005, 24'd7963435, 24'd8265005, 24'd8591036, 24'd8877007, 24'd9066325, 24'd9121523, 24'd9031679, 24'd8814572, 24'd8513168, 24'd8187113, 24'd7900934, 24'd7711264, 24'd7655640, 24'd7745068, 24'd7961852, 24'd8263090, 24'd8589167, 24'd8875555, 24'd9065576, 24'd9121626, 24'd9032614, 24'd8816153, 24'd8515083, 
24'd8188983, 24'd7902388, 24'd7712015, 24'd7655539, 24'd7744136, 24'd7960272, 24'd8261175, 24'd8587297, 24'd8874099, 24'd9064822, 24'd9121724, 24'd9033544, 24'd8817732, 24'd8516997, 24'd8190854, 24'd7903846, 24'd7712771, 24'd7655443, 24'd7743208, 24'd7958695, 24'd8259262, 24'd8585425, 24'd8872639, 24'd9064064, 24'd9121817, 24'd9034470, 24'd8819307, 24'd8518910, 24'd8192726, 24'd7905307, 
24'd7713532, 24'd7655353, 24'd7742284, 24'd7957121, 24'd8257349, 24'd8583552, 24'd8871176, 24'd9063301, 24'd9121905, 24'd9035391, 24'd8820879, 24'd8520822, 24'd8194600, 24'd7906771, 24'd7714297, 24'd7655268, 24'd7741365, 24'd7955551, 24'd8255437, 24'd8581678, 24'd8869710, 24'd9062533, 24'd9121988, 24'd9036308, 24'd8822449, 24'd8522733, 24'd8196475, 24'd7908239, 24'd7715067, 24'd7655188, 
24'd7740451, 24'd7953983, 24'd8253526, 24'd8579802, 24'd8868241, 24'd9061761, 24'd9122065, 24'd9037220, 24'd8824015, 24'd8524644, 24'd8198351, 24'd7909710, 24'd7715842, 24'd7655113, 24'd7739541, 24'd7952418, 24'd8251616, 24'd8577925, 24'd8866768, 24'd9060984, 24'd9122138, 24'd9038127, 24'd8825578, 24'd8526553, 24'd8200229, 24'd7911185, 24'd7716622, 24'd7655043, 24'd7738636, 24'd7950857, 
24'd8249707, 24'd8576046, 24'd8865292, 24'd9060202, 24'd9122205, 24'd9039030, 24'd8827138, 24'd8528462, 24'd8202108, 24'd7912663, 24'd7717406, 24'd7654979, 24'd7737735, 24'd7949298, 24'd8247799, 24'd8574167, 24'd8863812, 24'd9059415, 24'd9122267, 24'd9039929, 24'd8828695, 24'd8530369, 24'd8203989, 24'd7914144, 24'd7718195, 24'd7654919, 24'd7736839, 24'd7947742, 24'd8245892, 24'd8572285, 
24'd8862329, 24'd9058624, 24'd9122324, 24'd9040823, 24'd8830249, 24'd8532276, 24'd8205871, 24'd7915629, 24'd7718989, 24'd7654865, 24'd7735947, 24'd7946190, 24'd8243986, 24'd8570403, 24'd8860843, 24'd9057828, 24'd9122376, 24'd9041712, 24'd8831800, 24'd8534181, 24'd8207754, 24'd7917117, 24'd7719787, 24'd7654816, 24'd7735060, 24'd7944641, 24'd8242082, 24'd8568519, 24'd8859353, 24'd9057027, 
24'd9122422, 24'd9042597, 24'd8833348, 24'd8536086, 24'd8209638, 24'd7918608, 24'd7720590, 24'd7654771, 24'd7734178, 24'd7943095, 24'd8240178, 24'd8566635, 24'd8857860, 24'd9056222, 24'd9122464, 24'd9043477, 24'd8834892, 24'd8537989, 24'd8211523, 24'd7920102, 24'd7721398, 24'd7654733, 24'd7733300, 24'd7941552, 24'd8238275, 24'd8564748, 24'd8856364, 24'd9055412, 24'd9122500, 24'd9044352, 
24'd8836434, 24'd8539891, 24'd8213410, 24'd7921600, 24'd7722210, 24'd7654699, 24'd7732427, 24'd7940012, 24'd8236373, 24'd8562861, 24'd8854865, 24'd9054597, 24'd9122531, 24'd9045223, 24'd8837972, 24'd8541793, 24'd8215298, 24'd7923101, 24'd7723027, 24'd7654670, 24'd7731558, 24'd7938475, 24'd8234472, 24'd8560972, 24'd8853362, 24'd9053778, 24'd9122557, 24'd9046090, 24'd8839507, 24'd8543693, 
24'd8217187, 24'd7924606, 24'd7723849, 24'd7654647, 24'd7730694, 24'd7936941, 24'd8232572, 24'd8559083, 24'd8851856, 24'd9052953, 24'd9122578, 24'd9046951, 24'd8841039, 24'd8545592, 24'd8219078, 24'd7926113, 24'd7724675, 24'd7654628, 24'd7729835, 24'd7935411, 24'd8230674, 24'd8557191, 24'd8850347, 24'd9052125, 24'd9122594, 24'd9047808, 24'd8842568, 24'd8547490, 24'd8220969, 24'd7927624, 
24'd7725506, 24'd7654615, 24'd7728980, 24'd7933883, 24'd8228776, 24'd8555299, 24'd8848834, 24'd9051291, 24'd9122604, 24'd9048661, 24'd8844094, 24'd8549387, 24'd8222862, 24'd7929138, 24'd7726342, 24'd7654607, 24'd7728130, 24'd7932359, 24'd8226880, 24'd8553406, 24'd8847319, 24'd9050453, 24'd9122610, 24'd9049509, 24'd8845616, 24'd8551283, 24'd8224756, 24'd7930655, 24'd7727182, 24'd7654604, 
24'd7727284, 24'd7930839, 24'd8224985, 24'd8551511, 24'd8845800, 24'd9049611, 24'd9122610, 24'd9050352, 24'd8847136, 24'd8553178, 24'd8226651, 24'd7932176, 24'd7728027, 24'd7654607, 24'd7726443, 24'd7929321, 24'd8223091, 24'd8549616, 24'd8844278, 24'd9048763, 24'd9122605, 24'd9051191, 24'd8848652, 24'd8555071, 24'd8228548, 24'd7933700, 24'd7728877, 24'd7654614, 24'd7725607, 24'd7927806, 
24'd8221198, 24'd8547719, 24'd8842752, 24'd9047911, 24'd9122595, 24'd9052025, 24'd8850165, 24'd8556963, 24'd8230445, 24'd7935226, 24'd7729731, 24'd7654627, 24'd7724775, 24'd7926295, 24'd8219306, 24'd8545821, 24'd8841224, 24'd9047055, 24'd9122580, 24'd9052854, 24'd8851674, 24'd8558855, 24'd8232343, 24'd7936757, 24'd7730590, 24'd7654644, 24'd7723948, 24'd7924787, 24'd8217415, 24'd8543922, 
24'd8839692, 24'd9046194, 24'd9122560, 24'd9053678, 24'd8853181, 24'd8560745, 24'd8234243, 24'd7938290, 24'd7731454, 24'd7654667, 24'd7723126, 24'd7923282, 24'd8215526, 24'd8542022, 24'd8838157, 24'd9045328, 24'd9122535, 24'd9054498, 24'd8854684, 24'd8562633, 24'd8236144, 24'd7939826, 24'd7732322, 24'd7654695, 24'd7722308, 24'd7921781, 24'd8213638, 24'd8540121, 24'd8836619, 24'd9044457, 
24'd9122504, 24'd9055314, 24'd8856184, 24'd8564521, 24'd8238045, 24'd7941366, 24'd7733194, 24'd7654728, 24'd7721495, 24'd7920283, 24'd8211751, 24'd8538218, 24'd8835078, 24'd9043582, 24'd9122468, 24'd9056124, 24'd8857680, 24'd8566407, 24'd8239948, 24'd7942908, 24'd7734072, 24'd7654767, 24'd7720687, 24'd7918788, 24'd8209865, 24'd8536315, 24'd8833534, 24'd9042703, 24'd9122427, 24'd9056930, 
24'd8859173, 24'd8568292, 24'd8241852, 24'd7944454, 24'd7734954, 24'd7654810, 24'd7719883, 24'd7917296, 24'd8207981, 24'd8534411, 24'd8831987, 24'd9041819, 24'd9122381, 24'd9057732, 24'd8860663, 24'd8570176, 24'd8243757, 24'd7946003, 24'd7735840, 24'd7654859, 24'd7719085, 24'd7915808, 24'd8206097, 24'd8532505, 24'd8830436, 24'd9040930, 24'd9122330, 24'd9058528, 24'd8862150, 24'd8572059, 
24'd8245663, 24'd7947555, 24'd7736731, 24'd7654912, 24'd7718290, 24'd7914323, 24'd8204216, 24'd8530599, 24'd8828883, 24'd9040037, 24'd9122274, 24'd9059320, 24'd8863633, 24'd8573940, 24'd8247569, 24'd7949110, 24'd7737627, 24'd7654971, 24'd7717501, 24'd7912841, 24'd8202335, 24'd8528692, 24'd8827326, 24'd9039139, 24'd9122213, 24'd9060107, 24'd8865113, 24'd8575820, 24'd8249477, 24'd7950668, 
24'd7738527, 24'd7655035, 24'd7716716, 24'd7911363, 24'd8200456, 24'd8526783, 24'd8825766, 24'd9038236, 24'd9122146, 24'd9060890, 24'd8866590, 24'd8577698, 24'd8251386, 24'd7952230, 24'd7739432, 24'd7655104, 24'd7715936, 24'd7909888, 24'd8198578, 24'd8524874, 24'd8824203, 24'd9037329, 24'd9122074, 24'd9061667, 24'd8868063, 24'd8579576, 24'd8253296, 24'd7953794, 24'd7740341, 24'd7655179, 
24'd7715160, 24'd7908416, 24'd8196701, 24'd8522964, 24'd8822638, 24'd9036418, 24'd9121997, 24'd9062440, 24'd8869533, 24'd8581452, 24'd8255207, 24'd7955361, 24'd7741255, 24'd7655258, 24'd7714390, 24'd7906948, 24'd8194826, 24'd8521053, 24'd8821069, 24'd9035502, 24'd9121915, 24'd9063209, 24'd8871000, 24'd8583326, 24'd8257118, 24'd7956932, 24'd7742173, 24'd7655343, 24'd7713624, 24'd7905483, 
24'd8192952, 24'd8519140, 24'd8819497, 24'd9034581, 24'd9121828, 24'd9063972, 24'd8872463, 24'd8585200, 24'd8259031, 24'd7958505, 24'd7743096, 24'd7655432, 24'd7712863, 24'd7904022, 24'd8191079, 24'd8517227, 24'd8817922, 24'd9033656, 24'd9121736, 24'd9064731, 24'd8873923, 24'd8587072, 24'd8260944, 24'd7960082, 24'd7744023, 24'd7655527, 24'd7712106, 24'd7902563, 24'd8189208, 24'd8515313, 
24'd8816344, 24'd9032726, 24'd9121638, 24'd9065485, 24'd8875379, 24'd8588942, 24'd8262859, 24'd7961661, 24'd7744955, 24'd7655627, 24'd7711354, 24'd7901109, 24'd8187338, 24'd8513399, 24'd8814763, 24'd9031792, 24'd9121536, 24'd9066235, 24'd8876832, 24'd8590811, 24'd8264774, 24'd7963244, 24'd7745892, 24'd7655732, 24'd7710607, 24'd7899658, 24'd8185470, 24'd8511483, 24'd8813179, 24'd9030853, 
24'd9121428, 24'd9066979, 24'd8878282, 24'd8592679, 24'd8266690, 24'd7964829, 24'd7746833, 24'd7655843, 24'd7709865, 24'd7898210, 24'd8183603, 24'd8509566, 24'd8811592, 24'd9029910, 24'd9121315, 24'd9067719, 24'd8879728, 24'd8594545, 24'd8268607, 24'd7966417, 24'd7747778, 24'd7655958, 24'd7709128, 24'd7896765, 24'd8181737, 24'd8507649, 24'd8810002, 24'd9028962, 24'd9121197, 24'd9068454, 
24'd8881171, 24'd8596410, 24'd8270525, 24'd7968009, 24'd7748728, 24'd7656079, 24'd7708395, 24'd7895324, 24'd8179873, 24'd8505731, 24'd8808409, 24'd9028010, 24'd9121074, 24'd9069185, 24'd8882610, 24'd8598273, 24'd8272444, 24'd7969603, 24'd7749683, 24'd7656204, 24'd7707667, 24'd7893887, 24'd8178011, 24'd8503812, 24'd8806814, 24'd9027053, 24'd9120946, 24'd9069910, 24'd8884046, 24'd8600135, 
24'd8274363, 24'd7971200, 24'd7750642, 24'd7656335, 24'd7706944, 24'd7892453, 24'd8176150, 24'd8501892, 24'd8805215, 24'd9026092, 24'd9120813, 24'd9070631, 24'd8885478, 24'd8601995, 24'd8276284, 24'd7972801, 24'd7751605, 24'd7656471, 24'd7706226, 24'd7891022, 24'd8174290, 24'd8499971, 24'd8803613, 24'd9025127, 24'd9120674, 24'd9071347, 24'd8886907, 24'd8603854, 24'd8278205, 24'd7974404, 
24'd7752573, 24'd7656612, 24'd7705512, 24'd7889595, 24'd8172432, 24'd8498049, 24'd8802009, 24'd9024157, 24'd9120530, 24'd9072058, 24'd8888332, 24'd8605712, 24'd8280127, 24'd7976010, 24'd7753545, 24'd7656758, 24'd7704803, 24'd7888172, 24'd8170575, 24'd8496127, 24'd8800401, 24'd9023182, 24'd9120382, 24'd9072765, 24'd8889754, 24'd8607567, 24'd8282049, 24'd7977619, 24'd7754522, 24'd7656910, 
24'd7704099, 24'd7886751, 24'd8168720, 24'd8494204, 24'd8798791, 24'd9022203, 24'd9120228, 24'd9073466, 24'd8891172, 24'd8609422, 24'd8283973, 24'd7979230, 24'd7755503, 24'd7657066, 24'd7703400, 24'd7885335, 24'd8166867, 24'd8492281, 24'd8797178, 24'd9021220, 24'd9120069, 24'd9074163, 24'd8892587, 24'd8611275, 24'd8285897, 24'd7980845, 24'd7756489, 24'd7657228, 24'd7702705, 24'd7883922, 
24'd8165015, 24'd8490356, 24'd8795562, 24'd9020232, 24'd9119904, 24'd9074855, 24'd8893998, 24'd8613126, 24'd8287821, 24'd7982462, 24'd7757479, 24'd7657395, 24'd7702016, 24'd7882512, 24'd8163164, 24'd8488431, 24'd8793943, 24'd9019239, 24'd9119735, 24'd9075542, 24'd8895406, 24'd8614975, 24'd8289747, 24'd7984083, 24'd7758473, 24'd7657566, 24'd7701331, 24'd7881106, 24'd8161315, 24'd8486505, 
24'd8792321, 24'd9018243, 24'd9119561, 24'd9076225, 24'd8896810, 24'd8616823, 24'd8291673, 24'd7985706, 24'd7759472, 24'd7657743, 24'd7700651, 24'd7879704, 24'd8159468, 24'd8484578, 24'd8790696, 24'd9017242, 24'd9119381, 24'd9076902, 24'd8898211, 24'd8618670, 24'd8293600, 24'd7987332, 24'd7760476, 24'd7657926, 24'd7699976, 24'd7878305, 24'd8157623, 24'd8482651, 24'd8789069, 24'd9016236, 
24'd9119196, 24'd9077575, 24'd8899608, 24'd8620515, 24'd8295528, 24'd7988961, 24'd7761483, 24'd7658113, 24'd7699306, 24'd7876910, 24'd8155779, 24'd8480723, 24'd8787439, 24'd9015226, 24'd9119007, 24'd9078243, 24'd8901001, 24'd8622358, 24'd8297456, 24'd7990592, 24'd7762496, 24'd7658305, 24'd7698640, 24'd7875518, 24'd8153936, 24'd8478795, 24'd8785806, 24'd9014212, 24'd9118812, 24'd9078906, 
24'd8902391, 24'd8624199, 24'd8299385, 24'd7992227, 24'd7763512, 24'd7658503, 24'd7697979, 24'd7874130, 24'd8152095, 24'd8476866, 24'd8784170, 24'd9013193, 24'd9118612, 24'd9079564, 24'd8903777, 24'd8626039, 24'd8301314, 24'd7993864, 24'd7764533, 24'd7658705, 24'd7697324, 24'd7872746, 24'd8150256, 24'd8474936, 24'd8782531, 24'd9012170, 24'd9118407, 24'd9080217, 24'd8905160, 24'd8627878, 
24'd8303244, 24'd7995504, 24'd7765558, 24'd7658913, 24'd7696673, 24'd7871365, 24'd8148419, 24'd8473006, 24'd8780890, 24'd9011142, 24'd9118196, 24'd9080866, 24'd8906539, 24'd8629714, 24'd8305175, 24'd7997147, 24'd7766588, 24'd7659126, 24'd7696027, 24'd7869988, 24'd8146583, 24'd8471075, 24'd8779246, 24'd9010111, 24'd9117981, 24'd9081510, 24'd8907914, 24'd8631549, 24'd8307106, 24'd7998792, 
24'd7767622, 24'd7659344, 24'd7695385, 24'd7868614, 24'd8144749, 24'd8469143, 24'd8777599, 24'd9009074, 24'd9117760, 24'd9082148, 24'd8909286, 24'd8633382, 24'd8309038, 24'd8000440, 24'd7768660, 24'd7659567, 24'd7694749, 24'd7867245, 24'd8142917, 24'd8467211, 24'd8775949, 24'd9008034, 24'd9117535, 24'd9082782, 24'd8910654, 24'd8635214, 24'd8310970, 24'd8002091, 24'd7769703, 24'd7659795, 
24'd7694117, 24'd7865878, 24'd8141086, 24'd8465278, 24'd8774297, 24'd9006989, 24'd9117304, 24'd9083411, 24'd8912019, 24'd8637043, 24'd8312903, 24'd8003745, 24'd7770750, 24'd7660028, 24'd7693491, 24'd7864516, 24'd8139257, 24'd8463345, 24'd8772642, 24'd9005940, 24'd9117068, 24'd9084036, 24'd8913379, 24'd8638871, 24'd8314837, 24'd8005401, 24'd7771802, 24'd7660267, 24'd7692869, 24'd7863157, 
24'd8137430, 24'd8461411, 24'd8770984, 24'd9004886, 24'd9116827, 24'd9084655, 24'd8914736, 24'd8640698, 24'd8316771, 24'd8007060, 24'd7772857, 24'd7660510, 24'd7692252, 24'd7861802, 24'd8135605, 24'd8459477, 24'd8769324, 24'd9003828, 24'd9116581, 24'd9085270, 24'd8916090, 24'd8642522, 24'd8318705, 24'd8008722, 24'd7773917, 24'd7660759, 24'd7691640, 24'd7860450, 24'd8133781, 24'd8457542, 
24'd8767661, 24'd9002766, 24'd9116330, 24'd9085879, 24'd8917439, 24'd8644345, 24'd8320640, 24'd8010386, 24'd7774982, 24'd7661012, 24'd7691033, 24'd7859102, 24'd8131959, 24'd8455607, 24'd8765995, 24'd9001699, 24'd9116074, 24'd9086484, 24'd8918785, 24'd8646166, 24'd8322576, 24'd8012053, 24'd7776050, 24'd7661271, 24'd7690431, 24'd7857758, 24'd8130139, 24'd8453671, 24'd8764327, 24'd9000629, 
24'd9115812, 24'd9087084, 24'd8920128, 24'd8647985, 24'd8324512, 24'd8013723, 24'd7777123, 24'd7661535, 24'd7689833, 24'd7856418, 24'd8128321, 24'd8451735, 24'd8762656, 24'd8999554, 24'd9115546, 24'd9087678, 24'd8921466, 24'd8649802, 24'd8326448, 24'd8015395, 24'd7778201, 24'd7661804, 24'd7689241, 24'd7855081, 24'd8126505, 24'd8449799, 24'd8760983, 24'd8998474, 24'd9115274, 24'd9088268, 
24'd8922801, 24'd8651618, 24'd8328385, 24'd8017070, 24'd7779282, 24'd7662078, 24'd7688653, 24'd7853748, 24'd8124690, 24'd8447862, 24'd8759306, 24'd8997391, 24'd9114998, 24'd9088854, 24'd8924132, 24'd8653431, 24'd8330322, 24'd8018748, 24'd7780368, 24'd7662358, 24'd7688071, 24'd7852419, 24'd8122878, 24'd8445924, 24'd8757628, 24'd8996303, 24'd9114716, 24'd9089434, 24'd8925459, 24'd8655243, 
24'd8332260, 24'd8020428, 24'd7781458, 24'd7662642, 24'd7687493, 24'd7851093, 24'd8121067, 24'd8443986, 24'd8755946, 24'd8995210, 24'd9114429, 24'd9090009, 24'd8926783, 24'd8657053, 24'd8334198, 24'd8022110, 24'd7782552, 24'd7662931, 24'd7686920, 24'd7849772, 24'd8119258, 24'd8442048, 24'd8754262, 24'd8994114, 24'd9114137, 24'd9090579, 24'd8928103, 24'd8658861, 24'd8336136, 24'd8023796, 
24'd7783651, 24'd7663226, 24'd7686352, 24'd7848454, 24'd8117451, 24'd8440109, 24'd8752576, 24'd8993013, 24'd9113840, 24'd9091145, 24'd8929419, 24'd8660667, 24'd8338075, 24'd8025484, 24'd7784754, 24'd7663525, 24'd7685789, 24'd7847140, 24'd8115646, 24'd8438170, 24'd8750887, 24'd8991908, 24'd9113538, 24'd9091705, 24'd8930731, 24'd8662471, 24'd8340014, 24'd8027174, 24'd7785861, 24'd7663830, 
24'd7685231, 24'd7845830, 24'd8113843, 24'd8436231, 24'd8749195, 24'd8990799, 24'd9113231, 24'd9092261, 24'd8932039, 24'd8664273, 24'd8341954, 24'd8028867, 24'd7786972, 24'd7664140, 24'd7684678, 24'd7844523, 24'd8112041, 24'd8434291, 24'd8747501, 24'd8989686, 24'd9112919, 24'd9092812, 24'd8933344, 24'd8666074, 24'd8343893, 24'd8030562, 24'd7788087, 24'd7664454, 24'd7684130, 24'd7843220, 
24'd8110242, 24'd8432352, 24'd8745804, 24'd8988568, 24'd9112601, 24'd9093357, 24'd8934644, 24'd8667872, 24'd8345834, 24'd8032260, 24'd7789207, 24'd7664774, 24'd7683587, 24'd7841922, 24'd8108445, 24'd8430411, 24'd8744105, 24'd8987447, 24'd9112279, 24'd9093898, 24'd8935941, 24'd8669668, 24'd8347774, 24'd8033960, 24'd7790331, 24'd7665099, 24'd7683048, 24'd7840627, 24'd8106649, 24'd8428471, 
24'd8742403, 24'd8986321, 24'd9111951, 24'd9094434, 24'd8937234, 24'd8671463, 24'd8349715, 24'd8035663, 24'd7791459, 24'd7665429, 24'd7682515, 24'd7839335, 24'd8104856, 24'd8426530, 24'd8740699, 24'd8985190, 24'd9111619, 24'd9094965, 24'd8938524, 24'd8673255, 24'd8351656, 24'd8037369, 24'd7792591, 24'd7665764, 24'd7681987, 24'd7838048, 24'd8103064, 24'd8424589, 24'd8738993, 24'd8984056, 
24'd9111281, 24'd9095491, 24'd8939809, 24'd8675046, 24'd8353597, 24'd8039077, 24'd7793728, 24'd7666105, 24'd7681463, 24'd7836765, 24'd8101275, 24'd8422647, 24'd8737284, 24'd8982917, 24'd9110938, 24'd9096012, 24'd8941091, 24'd8676834, 24'd8355538, 24'd8040787, 24'd7794868, 24'd7666450, 24'd7680945, 24'd7835485, 24'd8099487, 24'd8420706, 24'd8735572, 24'd8981775, 24'd9110591, 24'd9096528, 
24'd8942368, 24'd8678621, 24'd8357480, 24'd8042500, 24'd7796013, 24'd7666800, 24'd7680431, 24'd7834209, 24'd8097702, 24'd8418764, 24'd8733858, 24'd8980628, 24'd9110238, 24'd9097039, 24'd8943642, 24'd8680405, 24'd8359422, 24'd8044215, 24'd7797162, 24'd7667155, 24'd7679923, 24'd7832938, 24'd8095918, 24'd8416822, 24'd8732142, 24'd8979477, 24'd9109880, 24'd9097545, 24'd8944912, 24'd8682188, 
24'd8361364, 24'd8045932, 24'd7798315, 24'd7667516, 24'd7679419, 24'd7831670, 24'd8094137, 24'd8414880, 24'd8730423, 24'd8978322, 24'd9109517, 24'd9098046, 24'd8946178, 24'd8683968, 24'd8363307, 24'd8047652, 24'd7799472, 24'd7667881, 24'd7678921, 24'd7830406, 24'd8092358, 24'd8412937, 24'd8728702, 24'd8977162, 24'd9109149, 24'd9098542, 24'd8947440, 24'd8685746, 24'd8365249, 24'd8049375, 
24'd7800634, 24'd7668252, 24'd7678427, 24'd7829146, 24'd8090581, 24'd8410995, 24'd8726978, 24'd8975999, 24'd9108776, 24'd9099033, 24'd8948698, 24'd8687522, 24'd8367192, 24'd8051099, 24'd7801799, 24'd7668627, 24'd7677938, 24'd7827889, 24'd8088805, 24'd8409052, 24'd8725252, 24'd8974831, 24'd9108398, 24'd9099519, 24'd8949952, 24'd8689296, 24'd8369135, 24'd8052826, 24'd7802969, 24'd7669008, 
24'd7677455, 24'd7826637, 24'd8087032, 24'd8407109, 24'd8723524, 24'd8973660, 24'd9108015, 24'd9100000, 24'd8951203, 24'd8691068, 24'd8371078, 24'd8054556, 24'd7804143, 24'd7669394, 24'd7676976, 24'd7825389, 24'd8085262, 24'd8405166, 24'd8721793, 24'd8972484, 24'd9107627, 24'd9100477, 24'd8952449, 24'd8692838, 24'd8373021, 24'd8056288, 24'd7805320, 24'd7669784, 24'd7676502, 24'd7824144, 
24'd8083493, 24'd8403223, 24'd8720061, 24'd8971304, 24'd9107233, 24'd9100948, 24'd8953691, 24'd8694606, 24'd8374964, 24'd8058022, 24'd7806502, 24'd7670180, 24'd7676034, 24'd7822904, 24'd8081726, 24'd8401280, 24'd8718325, 24'd8970120, 24'd9106835, 24'd9101414, 24'd8954930, 24'd8696371, 24'd8376907, 24'd8059758, 24'd7807688, 24'd7670581, 24'd7675570, 24'd7821668, 24'd8079962, 24'd8399336, 
24'd8716588, 24'd8968932, 24'd9106432, 24'd9101875, 24'd8956164, 24'd8698135, 24'd8378850, 24'd8061497, 24'd7808878, 24'd7670987, 24'd7675111, 24'd7820435, 24'd8078199, 24'd8397393, 24'd8714848, 24'd8967740, 24'd9106023, 24'd9102331, 24'd8957395, 24'd8699896, 24'd8380794, 24'd8063238, 24'd7810072, 24'd7671398, 24'd7674657, 24'd7819207, 24'd8076439, 24'd8395449, 24'd8713106, 24'd8966544, 
24'd9105610, 24'd9102783, 24'd8958621, 24'd8701655, 24'd8382737, 24'd8064981, 24'd7811270, 24'd7671813, 24'd7674209, 24'd7817982, 24'd8074681, 24'd8393506, 24'd8711361, 24'd8965344, 24'd9105192, 24'd9103229, 24'd8959844, 24'd8703412, 24'd8384681, 24'd8066727, 24'd7812473, 24'd7672234, 24'd7673765, 24'd7816762, 24'd8072926, 24'd8391562, 24'd8709614, 24'd8964140, 24'd9104768, 24'd9103670, 
24'd8961062, 24'd8705166, 24'd8386624, 24'd8068475, 24'd7813679, 24'd7672660, 24'd7673326, 24'd7815545, 24'd8071172, 24'd8389619, 24'd8707865, 24'd8962931, 24'd9104340, 24'd9104106, 24'd8962277, 24'd8706919, 24'd8388568, 24'd8070225, 24'd7814889, 24'd7673091, 24'd7672893, 24'd7814333, 24'd8069421, 24'd8387675, 24'd8706114, 24'd8961719, 24'd9103906, 24'd9104537, 24'd8963487, 24'd8708669, 
24'd8390512, 24'd8071977, 24'd7816104, 24'd7673527, 24'd7672464, 24'd7813124, 24'd8067672, 24'd8385732, 24'd8704361, 24'd8960503, 24'd9103468, 24'd9104963, 24'd8964693, 24'd8710417, 24'd8392455, 24'd8073732, 24'd7817322, 24'd7673968, 24'd7672040, 24'd7811920, 24'd8065925, 24'd8383788, 24'd8702605, 24'd8959282, 24'd9103024, 24'd9105385, 24'd8965896, 24'd8712163, 24'd8394399, 24'd8075489, 
24'd7818544, 24'd7674414, 24'd7671622, 24'd7810720, 24'd8064180, 24'd8381845, 24'd8700847, 24'd8958058, 24'd9102576, 24'd9105801, 24'd8967094, 24'd8713906, 24'd8396342, 24'd8077248, 24'd7819770, 24'd7674865, 24'd7671208, 24'd7809523, 24'd8062438, 24'd8379901, 24'd8699087, 24'd8956830, 24'd9102122, 24'd9106212, 24'd8968288, 24'd8715647, 24'd8398286, 24'd8079009, 24'd7821001, 24'd7675321, 
24'd7670800, 24'd7808331, 24'd8060698, 24'd8377958, 24'd8697325, 24'd8955598, 24'd9101664, 24'd9106618, 24'd8969479, 24'd8717386, 24'd8400229, 24'd8080772, 24'd7822235, 24'd7675782, 24'd7670396, 24'd7807143, 24'd8058960, 24'd8376014, 24'd8695561, 24'd8954361, 24'd9101200, 24'd9107019, 24'd8970665, 24'd8719123, 24'd8402172, 24'd8082537, 24'd7823473, 24'd7676248, 24'd7669998, 24'd7805959, 
24'd8057225, 24'd8374071, 24'd8693794, 24'd8953121, 24'd9100732, 24'd9107415, 24'd8971847, 24'd8720857, 24'd8404116, 24'd8084305, 24'd7824716, 24'd7676719, 24'd7669604, 24'd7804779, 24'd8055492, 24'd8372128, 24'd8692025, 24'd8951877, 24'd9100258, 24'd9107806, 24'd8973025, 24'd8722589, 24'd8406059, 24'd8086075, 24'd7825962, 24'd7677195, 24'd7669216, 24'd7803603, 24'd8053761, 24'd8370185, 
24'd8690254, 24'd8950629, 24'd9099780, 24'd9108191, 24'd8974199, 24'd8724318, 24'd8408002, 24'd8087847, 24'd7827212, 24'd7677676, 24'd7668833, 24'd7802431, 24'd8052033, 24'd8368242, 24'd8688482, 24'd8949377, 24'd9099296, 24'd9108572, 24'd8975368, 24'd8726046, 24'd8409944, 24'd8089621, 24'd7828466, 24'd7678162, 24'd7668454, 24'd7801263, 24'd8050307, 24'd8366299, 24'd8686707, 24'd8948121, 
24'd9098808, 24'd9108948, 24'd8976534, 24'd8727770, 24'd8411887, 24'd8091397, 24'd7829724, 24'd7678653, 24'd7668081, 24'd7800100, 24'd8048583, 24'd8364357, 24'd8684929, 24'd8946861, 24'd9098315, 24'd9109319, 24'd8977696, 24'd8729493, 24'd8413830, 24'd8093175, 24'd7830986, 24'd7679149, 24'd7667713, 24'd7798940, 24'd8046862, 24'd8362414, 24'd8683150, 24'd8945597, 24'd9097816, 24'd9109684, 
24'd8978853, 24'd8731213, 24'd8415772, 24'd8094955, 24'd7832252, 24'd7679650, 24'd7667350, 24'd7797785, 24'd8045143, 24'd8360472, 24'd8681369, 24'd8944329, 24'd9097313, 24'd9110045, 24'd8980006, 24'd8732931, 24'd8417714, 24'd8096737, 24'd7833521, 24'd7680156, 24'd7666992, 24'd7796634, 24'd8043426, 24'd8358530, 24'd8679586, 24'd8943057, 24'd9096804, 24'd9110401, 24'd8981155, 24'd8734646, 
24'd8419656, 24'd8098522, 24'd7834795, 24'd7680667, 24'd7666638, 24'd7795487, 24'd8041712, 24'd8356588, 24'd8677800, 24'd8941782, 24'd9096291, 24'd9110751, 24'd8982300, 24'd8736359, 24'd8421598, 24'd8100308, 24'd7836072, 24'd7681182, 24'd7666291, 24'd7794344, 24'd8040001, 24'd8354646, 24'd8676013, 24'd8940502, 24'd9095773, 24'd9111097, 24'd8983441, 24'd8738069, 24'd8423539, 24'd8102097, 
24'd7837354, 24'd7681703, 24'd7665948, 24'd7793205, 24'd8038292, 24'd8352705, 24'd8674224, 24'd8939219, 24'd9095250, 24'd9111437, 24'd8984578, 24'd8739777, 24'd8425480, 24'd8103887, 24'd7838639, 24'd7682229, 24'd7665610, 24'd7792071, 24'd8036585, 24'd8350764, 24'd8672432, 24'd8937932, 24'd9094721, 24'd9111772, 24'd8985710, 24'd8741482, 24'd8427421, 24'd8105679, 24'd7839928, 24'd7682760, 
24'd7665277, 24'd7790940, 24'd8034881, 24'd8348823, 24'd8670639, 24'd8936641, 24'd9094188, 24'd9112102, 24'd8986838, 24'd8743185, 24'd8429362, 24'd8107474, 24'd7841221, 24'd7683295, 24'd7664949, 24'd7789814, 24'd8033179, 24'd8346883, 24'd8668843, 24'd8935346, 24'd9093650, 24'd9112428, 24'd8987962, 24'd8744886, 24'd8431303, 24'd8109270, 24'd7842518, 24'd7683836, 24'd7664627, 24'd7788692, 
24'd8031480, 24'd8344942, 24'd8667046, 24'd8934047, 24'd9093107, 24'd9112748, 24'd8989082, 24'd8746584, 24'd8433243, 24'd8111068, 24'd7843818, 24'd7684381, 24'd7664309, 24'd7787574, 24'd8029783, 24'd8343002, 24'd8665247, 24'd8932745, 24'd9092559, 24'd9113063, 24'd8990198, 24'd8748279, 24'd8435183, 24'd8112869, 24'd7845123, 24'd7684932, 24'd7663997, 24'd7786461, 24'd8028089, 24'd8341063, 
24'd8663446, 24'd8931439, 24'd9092006, 24'd9113373, 24'd8991309, 24'd8749972, 24'd8437122, 24'd8114671, 24'd7846431, 24'd7685487, 24'd7663689, 24'd7785352, 24'd8026397, 24'd8339123, 24'd8661642, 24'd8930128, 24'd9091448, 24'd9113677, 24'd8992417, 24'd8751663, 24'd8439061, 24'd8116475, 24'd7847743, 24'd7686047, 24'd7663387, 24'd7784246, 24'd8024708, 24'd8337184, 24'd8659837, 24'd8928814, 
24'd9090886, 24'd9113977, 24'd8993520, 24'd8753351, 24'd8441000, 24'd8118281, 24'd7849059, 24'd7686613, 24'd7663090, 24'd7783146, 24'd8023021, 24'd8335246, 24'd8658030, 24'd8927497, 24'd9090318, 24'd9114272, 24'd8994618, 24'd8755036, 24'd8442938, 24'd8120089, 24'd7850379, 24'd7687183, 24'd7662798, 24'd7782049, 24'd8021337, 24'd8333307, 24'd8656222, 24'd8926175, 24'd9089745, 24'd9114562, 
24'd8995713, 24'd8756719, 24'd8444877, 24'd8121899, 24'd7851702, 24'd7687758, 24'd7662511, 24'd7780957, 24'd8019656, 24'd8331370, 24'd8654411, 24'd8924850, 24'd9089168, 24'd9114846, 24'd8996803, 24'd8758399, 24'd8446814, 24'd8123710, 24'd7853029, 24'd7688338, 24'd7662229, 24'd7779869, 24'd8017977, 24'd8329432, 24'd8652598, 24'd8923521, 24'd9088585, 24'd9115125, 24'd8997889, 24'd8760077, 
24'd8448751, 24'd8125524, 24'd7854360, 24'd7688923, 24'd7661952, 24'd7778785, 24'd8016300, 24'd8327495, 24'd8650784, 24'd8922188, 24'd9087998, 24'd9115400, 24'd8998971, 24'd8761752, 24'd8450688, 24'd8127339, 24'd7855695, 24'd7689512, 24'd7661680, 24'd7777705, 24'd8014627, 24'd8325558, 24'd8648967, 24'd8920852, 24'd9087406, 24'd9115669, 24'd9000048, 24'd8763424, 24'd8452625, 24'd8129156, 
24'd7857033, 24'd7690107, 24'd7661413, 24'd7776630, 24'd8012956, 24'd8323622, 24'd8647149, 24'd8919511, 24'd9086809, 24'd9115933, 24'd9001121, 24'd8765094, 24'd8454561, 24'd8130975, 24'd7858375, 24'd7690707, 24'd7661152, 24'd7775559, 24'd8011287, 24'd8321687, 24'd8645329, 24'd8918167, 24'd9086207, 24'd9116192, 24'd9002190, 24'd8766761, 24'd8456496, 24'd8132796, 24'd7859721, 24'd7691311, 
24'd7660895, 24'd7774492, 24'd8009621, 24'd8319751, 24'd8643508, 24'd8916820, 24'd9085600, 24'd9116446, 24'd9003254, 24'd8768425, 24'd8458431, 24'd8134619, 24'd7861070, 24'd7691921, 24'd7660644, 24'd7773430, 24'd8007958, 24'd8317817, 24'd8641684, 24'd8915468, 24'd9084988, 24'd9116695, 24'd9004315, 24'd8770087, 24'd8460366, 24'd8136443, 24'd7862424, 24'd7692535, 24'd7660398, 24'd7772372, 
24'd8006298, 24'd8315882, 24'd8639859, 24'd8914113, 24'd9084371, 24'd9116939, 24'd9005371, 24'd8771746, 24'd8462300, 24'd8138269, 24'd7863781, 24'd7693154, 24'd7660157, 24'd7771318, 24'd8004640, 24'd8313949, 24'd8638032, 24'd8912755, 24'd9083750, 24'd9117177, 24'd9006422, 24'd8773403, 24'd8464233, 24'd8140097, 24'd7865141, 24'd7693778, 24'd7659920, 24'd7770269, 24'd8002985, 24'd8312015, 
24'd8636203, 24'd8911392, 24'd9083123, 24'd9117411, 24'd9007469, 24'd8775057, 24'd8466166, 24'd8141927, 24'd7866505, 24'd7694407, 24'd7659690, 24'd7769224, 24'd8001333, 24'd8310083, 24'd8634373, 24'd8910026, 24'd9082492, 24'd9117639, 24'd9008512, 24'd8776708, 24'd8468099, 24'd8143758, 24'd7867873, 24'd7695041, 24'd7659464, 24'd7768183, 24'd7999683, 24'd8308150, 24'd8632540, 24'd8908656, 
24'd9081856, 24'd9117862, 24'd9009551, 24'd8778356, 24'd8470030, 24'd8145591, 24'd7869245, 24'd7695679, 24'd7659243, 24'd7767146, 24'd7998036, 24'd8306219, 24'd8630706, 24'd8907283, 24'd9081215, 24'd9118080, 24'd9010585, 24'd8780001, 24'd8471962, 24'd8147426, 24'd7870620, 24'd7696323, 24'd7659027, 24'd7766114, 24'd7996392, 24'd8304288, 24'd8628871, 24'd8905906, 24'd9080569, 24'd9118294, 
24'd9011615, 24'd8781644, 24'd8473892, 24'd8149263, 24'd7871999, 24'd7696971, 24'd7658817, 24'd7765087, 24'd7994750, 24'd8302357, 24'd8627033, 24'd8904525, 24'd9079918, 24'd9118501, 24'd9012640, 24'd8783284, 24'd8475823, 24'd8151101, 24'd7873382, 24'd7697624, 24'd7658612, 24'd7764064, 24'd7993112, 24'd8300428, 24'd8625194, 24'd8903141, 24'd9079262, 24'd9118704, 24'd9013661, 24'd8784922, 
24'd8477752, 24'd8152941, 24'd7874768, 24'd7698282, 24'd7658411, 24'd7763045, 24'd7991476, 24'd8298498, 24'd8623354, 24'd8901753, 24'd9078602, 24'd9118902, 24'd9014678, 24'd8786556, 24'd8479681, 24'd8154782, 24'd7876157, 24'd7698945, 24'd7658216, 24'd7762030, 24'd7989843, 24'd8296570, 24'd8621511, 24'd8900361, 24'd9077936, 24'd9119095, 24'd9015691, 24'd8788188, 24'd8481609, 24'd8156625, 
24'd7877551, 24'd7699613, 24'd7658026, 24'd7761020, 24'd7988212, 24'd8294642, 24'd8619667, 24'd8898966, 24'd9077266, 24'd9119282, 24'd9016698, 24'd8789817, 24'd8483537, 24'd8158470, 24'd7878947, 24'd7700286, 24'd7657841, 24'd7760014, 24'd7986585, 24'd8292715, 24'd8617822, 24'd8897568, 24'd9076591, 24'd9119464, 24'd9017702, 24'd8791443, 24'd8485464, 24'd8160317, 24'd7880348, 24'd7700963, 
24'd7657661, 24'd7759013, 24'd7984960, 24'd8290788, 24'd8615975, 24'd8896166, 24'd9075912, 24'd9119642, 24'd9018701, 24'd8793066, 24'd8487390, 24'd8162165, 24'd7881752, 24'd7701645, 24'd7657487, 24'd7758016, 24'd7983338, 24'd8288862, 24'd8614126, 24'd8894760, 24'd9075227, 24'd9119814, 24'd9019696, 24'd8794687, 24'd8489315, 24'd8164014, 24'd7883159, 24'd7702332, 24'd7657317, 24'd7757024, 
24'd7981719, 24'd8286937, 24'd8612275, 24'd8893350, 24'd9074538, 24'd9119981, 24'd9020686, 24'd8796304, 24'd8491240, 24'd8165865, 24'd7884571, 24'd7703024, 24'd7657153, 24'd7756035, 24'd7980103, 24'd8285013, 24'd8610424, 24'd8891938, 24'd9073843, 24'd9120142, 24'd9021672, 24'd8797919, 24'd8493164, 24'd8167718, 24'd7885985, 24'd7703720, 24'd7656994, 24'd7755052, 24'd7978490, 24'd8283089, 
24'd8608570, 24'd8890521, 24'd9073144, 24'd9120299, 24'd9022653, 24'd8799531, 24'd8495088, 24'd8169572, 24'd7887403, 24'd7704422, 24'd7656840, 24'd7754073, 24'd7976879, 24'd8281166, 24'd8606715, 24'd8889101, 24'd9072441, 24'd9120451, 24'd9023630, 24'd8801140, 24'd8497010, 24'd8171428, 24'd7888825, 24'd7705128, 24'd7656691, 24'd7753098, 24'd7975272, 24'd8279244, 24'd8604859, 24'd8887678, 
24'd9071732, 24'd9120597, 24'd9024603, 24'd8802746, 24'd8498932, 24'd8173285, 24'd7890250, 24'd7705839, 24'd7656547, 24'd7752128, 24'd7973667, 24'd8277322, 24'd8603000, 24'd8886251, 24'd9071019, 24'd9120738, 24'd9025571, 24'd8804349, 24'd8500853, 24'd8175144, 24'd7891679, 24'd7706555, 24'd7656408, 24'd7751162, 24'd7972065, 24'd8275401, 24'd8601141, 24'd8884820, 24'd9070300, 24'd9120875, 
24'd9026534, 24'd8805950, 24'd8502774, 24'd8177004, 24'd7893111, 24'd7707276, 24'd7656274, 24'd7750201, 24'd7970466, 24'd8273481, 24'd8599280, 24'd8883387, 24'd9069577, 24'd9121006, 24'd9027493, 24'd8807547, 24'd8504693, 24'd8178866, 24'd7894547, 24'd7708001, 24'd7656146, 24'd7749244, 24'd7968870, 24'd8271562, 24'd8597417, 24'd8881949, 24'd9068850, 24'd9121131, 24'd9028448, 24'd8809141, 
24'd8506612, 24'd8180730, 24'd7895986, 24'd7708731, 24'd7656023, 24'd7748291, 24'd7967277, 24'd8269644, 24'd8595553, 24'd8880508, 24'd9068117, 24'd9121252, 24'd9029398, 24'd8810733, 24'd8508530, 24'd8182594, 24'd7897428, 24'd7709466, 24'd7655904, 24'd7747343, 24'd7965687, 24'd8267727, 24'd8593688, 24'd8879064, 24'd9067380, 24'd9121368, 24'd9030344, 24'd8812321, 24'd8510447, 24'd8184460, 
24'd7898874, 24'd7710206, 24'd7655791, 24'd7746400, 24'd7964100, 24'd8265810, 24'd8591821, 24'd8877616, 24'd9066638, 24'd9121478, 24'd9031285, 24'd8813907, 24'd8512363, 24'd8186328, 24'd7900324, 24'd7710950, 24'd7655683, 24'd7745461, 24'd7962516, 24'd8263894, 24'd8589953, 24'd8876165, 24'd9065891, 24'd9121584, 24'd9032222, 24'd8815490, 24'd8514278, 24'd8188197, 24'd7901777, 24'd7711699, 
24'd7655581, 24'd7744527, 24'd7960935, 24'd8261979, 24'd8588083, 24'd8874711, 24'd9065139, 24'd9121684, 24'd9033154, 24'd8817069, 24'd8516193, 24'd8190068, 24'd7903233, 24'd7712453, 24'd7655483, 24'd7743597, 24'd7959357, 24'd8260065, 24'd8586212, 24'd8873253, 24'd9064383, 24'd9121779, 24'd9034081, 24'd8818646, 24'd8518106, 24'd8191939, 24'd7904693, 24'd7713212, 24'd7655390, 24'd7742671, 
24'd7957782, 24'd8258152, 24'd8584339, 24'd8871791, 24'd9063622, 24'd9121869, 24'd9035005, 24'd8820219, 24'd8520019, 24'd8193813, 24'd7906156, 24'd7713975, 24'd7655303, 24'd7741751, 24'd7956210, 24'd8256240, 24'd8582465, 24'd8870327, 24'd9062856, 24'd9121954, 24'd9035923, 24'd8821790, 24'd8521931, 24'd8195687, 24'd7907622, 24'd7714743, 24'd7655221, 24'd7740834, 24'd7954641, 24'd8254329, 
24'd8580590, 24'd8868858, 24'd9062086, 24'd9122033, 24'd9036837, 24'd8823357, 24'd8523841, 24'd8197563, 24'd7909092, 24'd7715516, 24'd7655144, 24'd7739923, 24'd7953075, 24'd8252418, 24'd8578714, 24'd8867387, 24'd9061311, 24'd9122108, 24'd9037747, 24'd8824922, 24'd8525751, 24'd8199440, 24'd7910565, 24'd7716294, 24'd7655072, 24'd7739015, 24'd7951512, 24'd8250509, 24'd8576836, 24'd8865912, 
24'd9060531, 24'd9122177, 24'd9038651, 24'd8826483, 24'd8527660, 24'd8201319, 24'd7912042, 24'd7717076, 24'd7655005, 24'd7738113, 24'd7949952, 24'd8248601, 24'd8574956, 24'd8864434, 24'd9059746, 24'd9122241, 24'd9039552, 24'd8828042, 24'd8529568, 24'd8203199, 24'd7913521, 24'd7717863, 24'd7654943, 24'd7737215, 24'd7948395, 24'd8246693, 24'd8573076, 24'd8862952, 24'd9058957, 24'd9122300, 
24'd9040448, 24'd8829597, 24'd8531475, 24'd8205080, 24'd7915005, 24'd7718655, 24'd7654887, 24'd7736321, 24'd7946842, 24'd8244787, 24'd8571194, 24'd8861467, 24'd9058163, 24'd9122354, 24'd9041339, 24'd8831149, 24'd8533381, 24'd8206962, 24'd7916491, 24'd7719451, 24'd7654836, 24'd7735432, 24'd7945291, 24'd8242882, 24'd8569311, 24'd8859979, 24'd9057364, 24'd9122403, 24'd9042225, 24'd8832698, 
24'd8535286, 24'd8208846, 24'd7917981, 24'd7720252, 24'd7654789, 24'd7734548, 24'd7943744, 24'd8240977, 24'd8567426, 24'd8858488, 24'd9056561, 24'd9122447, 24'd9043108, 24'd8834244, 24'd8537190, 24'd8210731, 24'd7919474, 24'd7721058, 24'd7654748, 24'd7733668, 24'd7942199, 24'd8239074, 24'd8565541, 24'd8856993, 24'd9055753, 24'd9122485, 24'd9043985, 24'd8835787, 24'd8539092, 24'd8212617, 
24'd7920971, 24'd7721868, 24'd7654712, 24'd7732793, 24'd7940658, 24'd8237172, 24'd8563654, 24'd8855495, 24'd9054940, 24'd9122519, 24'd9044858, 24'd8837326, 24'd8540994, 24'd8214505, 24'd7922470, 24'd7722683, 24'd7654682, 24'd7731922, 24'd7939120, 24'd8235270, 24'd8561766, 24'd8853994, 24'd9054122, 24'd9122547, 24'd9045726, 24'd8838863, 24'd8542895, 24'd8216394, 24'd7923973, 24'd7723503, 
24'd7654656, 24'd7731056, 24'd7937585, 24'd8233370, 24'd8559876, 24'd8852489, 24'd9053300, 24'd9122570, 24'd9046590, 24'd8840396, 24'd8544794, 24'd8218284, 24'd7925480, 24'd7724328, 24'd7654635, 24'd7730195, 24'd7936053, 24'd8231471, 24'd8557986, 24'd8850981, 24'd9052473, 24'd9122588, 24'd9047449, 24'd8841926, 24'd8546693, 24'd8220175, 24'd7926989, 24'd7725157, 24'd7654620, 24'd7729338, 
24'd7934525, 24'd8229573, 24'd8556094, 24'd8849470, 24'd9051642, 24'd9122601, 24'd9048303, 24'd8843453, 24'd8548590, 24'd8222067, 24'd7928502, 24'd7725990, 24'd7654610, 24'd7728486, 24'd7932999, 24'd8227676, 24'd8554201, 24'd8847956, 24'd9050806, 24'd9122608, 24'd9049153, 24'd8844977, 24'd8550487, 24'd8223961, 24'd7930018, 24'd7726829, 24'd7654605, 24'd7727639, 24'd7931477, 24'd8225781, 
24'd8552307, 24'd8846438, 24'd9049965, 24'd9122611, 24'd9049998, 24'd8846498, 24'd8552382, 24'd8225855, 24'd7931537, 24'd7727672, 24'd7654605, 24'd7726796, 24'd7929958, 24'd8223886, 24'd8550412, 24'd8844917, 24'd9049120, 24'd9122608, 24'd9050839, 24'd8848015, 24'd8554276, 24'd8227751, 24'd7933059, 24'd7728520, 24'd7654610, 24'd7725958, 24'd7928442, 24'd8221993, 24'd8548516, 24'd8843393, 
24'd9048270, 24'd9122600, 24'd9051675, 24'd8849530, 24'd8556169, 24'd8229648, 24'd7934585, 24'd7729372, 24'd7654621, 24'd7725124, 24'd7926930, 24'd8220100, 24'd8546618, 24'd8841866, 24'd9047415, 24'd9122587, 24'd9052506, 24'd8851041, 24'd8558060, 24'd8231546, 24'd7936113, 24'd7730229, 24'd7654636, 24'd7724295, 24'd7925420, 24'd8218209, 24'd8544720, 24'd8840336, 24'd9046556, 24'd9122569, 
24'd9053333, 24'd8852548, 24'd8559951, 24'd8233445, 24'd7937645, 24'd7731090, 24'd7654657, 24'd7723471, 24'd7923914, 24'd8216319, 24'd8542820, 24'd8838802, 24'd9045692, 24'd9122546, 24'd9054155, 24'd8854053, 24'd8561840, 24'd8235345, 24'd7939180, 24'd7731957, 24'd7654683, 24'd7722651, 24'd7922411, 24'd8214431, 24'd8540919, 24'd8837266, 24'd9044824, 24'd9122517, 24'd9054972, 24'd8855554, 
24'd8563728, 24'd8237246, 24'd7940719, 24'd7732827, 24'd7654714, 24'd7721836, 24'd7920912, 24'd8212543, 24'd8539018, 24'd8835726, 24'd9043951, 24'd9122484, 24'd9055784, 24'd8857052, 24'd8565615, 24'd8239149, 24'd7942260, 24'd7733703, 24'd7654750, 24'd7721026, 24'd7919415, 24'd8210657, 24'd8537115, 24'd8834183, 24'd9043073, 24'd9122445, 24'd9056592, 24'd8858547, 24'd8567501, 24'd8241052, 
24'd7943805, 24'd7734583, 24'd7654791, 24'd7720220, 24'd7917922, 24'd8208772, 24'd8535211, 24'd8832637, 24'd9042191, 24'd9122401, 24'd9057396, 24'd8860038, 24'd8569385, 24'd8242957, 24'd7945352, 24'd7735467, 24'd7654837, 24'd7719420, 24'd7916433, 24'd8206888, 24'd8533306, 24'd8831088, 24'd9041304, 24'd9122352, 24'd9058194, 24'd8861526, 24'd8571268, 24'd8244862, 24'd7946903, 24'd7736356, 
24'd7654889, 24'd7718623, 24'd7914946, 24'd8205006, 24'd8531400, 24'd8829536, 24'd9040412, 24'd9122298, 24'd9058988, 24'd8863011, 24'd8573150, 24'd8246768, 24'd7948457, 24'd7737250, 24'd7654946, 24'd7717832, 24'd7913463, 24'd8203125, 24'd8529493, 24'd8827980, 24'd9039516, 24'd9122239, 24'd9059777, 24'd8864492, 24'd8575030, 24'd8248676, 24'd7950014, 24'd7738148, 24'd7655008, 24'd7717045, 
24'd7911983, 24'd8201245, 24'd8527585, 24'd8826422, 24'd9038616, 24'd9122175, 24'd9060562, 24'd8865970, 24'd8576910, 24'd8250584, 24'd7951574, 24'd7739051, 24'd7655075, 24'd7716263, 24'd7910507, 24'd8199366, 24'd8525676, 24'd8824860, 24'd9037711, 24'd9122105, 24'd9061341, 24'd8867445, 24'd8578787, 24'd8252494, 24'd7953137, 24'd7739958, 24'd7655147, 24'd7715486, 24'd7909034, 24'd8197489, 
24'd8523766, 24'd8823296, 24'd9036801, 24'd9122030, 24'd9062116, 24'd8868916, 24'd8580664, 24'd8254404, 24'd7954703, 24'd7740870, 24'd7655224, 24'd7714713, 24'd7907564, 24'd8195613, 24'd8521855, 24'd8821728, 24'd9035887, 24'd9121950, 24'd9062887, 24'd8870384, 24'd8582539, 24'd8256315, 24'd7956272, 24'd7741787, 24'd7655306, 24'd7713945, 24'd7906098, 24'd8193739, 24'd8519944, 24'd8820157, 
24'd9034968, 24'd9121865, 24'd9063652, 24'd8871849, 24'd8584413, 24'd8258227, 24'd7957844, 24'd7742708, 24'd7655394, 24'd7713182, 24'd7904635, 24'd8191866, 24'd8518031, 24'd8818584, 24'd9034045, 24'd9121775, 24'd9064413, 24'd8873310, 24'd8586285, 24'd8260141, 24'd7959419, 24'd7743633, 24'd7655487, 24'd7712423, 24'd7903176, 24'd8189994, 24'd8516117, 24'd8817007, 24'd9033117, 24'd9121680, 
24'd9065169, 24'd8874768, 24'd8588156, 24'd8262055, 24'd7960997, 24'd7744563, 24'd7655585, 24'd7711670, 24'd7901719, 24'd8188124, 24'd8514203, 24'd8815427, 24'd9032185, 24'd9121580, 24'd9065921, 24'd8876222, 24'd8590026, 24'd8263970, 24'd7962579, 24'd7745498, 24'd7655688, 24'd7710921, 24'd7900267, 24'd8186255, 24'd8512288, 24'd8813845, 24'd9031248, 24'd9121474, 24'd9066667, 24'd8877673, 
24'd8591894, 24'd8265885, 24'd7964163, 24'd7746437, 24'd7655796, 24'd7710176, 24'd7898817, 24'd8184387, 24'd8510371, 24'd8812259, 24'd9030307, 24'd9121363, 24'd9067409, 24'd8879121, 24'd8593761, 24'd8267802, 24'd7965750, 24'd7747381, 24'd7655909, 24'd7709437, 24'd7897372, 24'd8182521, 24'd8508454, 24'd8810670, 24'd9029361, 24'd9121248, 24'd9068146, 24'd8880565, 24'd8595627, 24'd8269719, 
24'd7967340, 24'd7748329, 24'd7656027, 24'd7708702, 24'd7895929, 24'd8180656, 24'd8506536, 24'd8809079, 24'd9028411, 24'd9121127, 24'd9068878, 24'd8882006, 24'd8597491, 24'd8271638, 24'd7968933, 24'd7749281, 24'd7656151, 24'd7707972, 24'd7894490, 24'd8178793, 24'd8504618, 24'd8807484, 24'd9027456, 24'd9121000, 24'd9069606, 24'd8883443, 24'd8599353, 24'd8273557, 24'd7970529, 24'd7750238, 
24'd7656279, 24'd7707247, 24'd7893055, 24'd8176931, 24'd8502698, 24'd8805887, 24'd9026497, 24'd9120869, 24'd9070329, 24'd8884877, 24'd8601214, 24'd8275477, 24'd7972128, 24'd7751200, 24'd7656413, 24'd7706527, 24'd7891623, 24'd8175071, 24'd8500778, 24'd8804286, 24'd9025533, 24'd9120733, 24'd9071047, 24'd8886307, 24'd8603074, 24'd8277398, 24'd7973730, 24'd7752166, 24'd7656552, 24'd7705811, 
24'd7890194, 24'd8173212, 24'd8498857, 24'd8802683, 24'd9024565, 24'd9120591, 24'd9071760, 24'd8887734, 24'd8604932, 24'd8279319, 24'd7975335, 24'd7753136, 24'd7656696, 24'd7705100, 24'd7888769, 24'd8171355, 24'd8496935, 24'd8801077, 24'd9023592, 24'd9120445, 24'd9072468, 24'd8889157, 24'd8606788, 24'd8281241, 24'd7976942, 24'd7754111, 24'd7656845, 24'd7704394, 24'd7887348, 24'd8169499, 
24'd8495012, 24'd8799468, 24'd9022615, 24'd9120293, 24'd9073172, 24'd8890577, 24'd8608643, 24'd8283165, 24'd7978553, 24'd7755090, 24'd7657000, 24'd7703693, 24'd7885929, 24'd8167645, 24'd8493089, 24'd8797856, 24'd9021633, 24'd9120136, 24'd9073871, 24'd8891993, 24'd8610496, 24'd8285088, 24'd7980166, 24'd7756074, 24'd7657159, 24'd7702997, 24'd7884515, 24'd8165792, 24'd8491165, 24'd8796241, 
24'd9020647, 24'd9119974, 24'd9074565, 24'd8893406, 24'd8612348, 24'd8287013, 24'd7981783, 24'd7757062, 24'd7657324, 24'd7702305, 24'd7883104, 24'd8163941, 24'd8489240, 24'd8794623, 24'd9019657, 24'd9119807, 24'd9075254, 24'd8894815, 24'd8614199, 24'd8288938, 24'd7983402, 24'd7758055, 24'd7657494, 24'd7701618, 24'd7881697, 24'd8162092, 24'd8487314, 24'd8793002, 24'd9018662, 24'd9119635, 
24'd9075938, 24'd8896221, 24'd8616047, 24'd8290864, 24'd7985024, 24'd7759052, 24'd7657668, 24'd7700936, 24'd7880293, 24'd8160244, 24'd8485388, 24'd8791379, 24'd9017663, 24'd9119457, 24'd9076618, 24'd8897623, 24'd8617894, 24'd8292791, 24'd7986649, 24'd7760054, 24'd7657848, 24'd7700259, 24'd7878892, 24'd8158398, 24'd8483461, 24'd8789753, 24'd9016659, 24'd9119275, 24'd9077293, 24'd8899021, 
24'd8619740, 24'd8294718, 24'd7988276, 24'd7761060, 24'd7658033, 24'd7699587, 24'd7877496, 24'd8156553, 24'd8481533, 24'd8788124, 24'd9015651, 24'd9119087, 24'd9077963, 24'd8900416, 24'd8621584, 24'd8296646, 24'd7989907, 24'd7762070, 24'd7658224, 24'd7698919, 24'd7876103, 24'd8154710, 24'd8479605, 24'd8786492, 24'd9014638, 24'd9118894, 24'd9078628, 24'd8901808, 24'd8623426, 24'd8298574, 
24'd7991540, 24'd7763085, 24'd7658419, 24'd7698256, 24'd7874713, 24'd8152868, 24'd8477676, 24'd8784857, 24'd9013621, 24'd9118696, 24'd9079288, 24'd8903195, 24'd8625267, 24'd8300504, 24'd7993176, 24'd7764104, 24'd7658619, 24'd7697599, 24'd7873327, 24'd8151029, 24'd8475747, 24'd8783220, 24'd9012600, 24'd9118493, 24'd9079944, 24'd8904580, 24'd8627106, 24'd8302433, 24'd7994815, 24'd7765127, 
24'd7658825, 24'd7696946, 24'd7871945, 24'd8149190, 24'd8473816, 24'd8781580, 24'd9011574, 24'd9118285, 24'd9080594, 24'd8905960, 24'd8628943, 24'd8304364, 24'd7996456, 24'd7766155, 24'd7659036, 24'd7696297, 24'd7870566, 24'd8147354, 24'd8471886, 24'd8779937, 24'd9010544, 24'd9118072, 24'd9081240, 24'd8907337, 24'd8630779, 24'd8306295, 24'd7998101, 24'd7767187, 24'd7659252, 24'd7695654, 
24'd7869191, 24'd8145519, 24'd8469954, 24'd8778291, 24'd9009510, 24'd9117854, 24'd9081881, 24'd8908710, 24'd8632612, 24'd8308226, 24'd7999748, 24'd7768224, 24'd7659472, 24'd7695016, 24'd7867819, 24'd8143686, 24'd8468022, 24'd8776643, 24'd9008471, 24'd9117630, 24'd9082517, 24'd8910080, 24'd8634445, 24'd8310159, 24'd8001398, 24'd7769265, 24'd7659699, 24'd7694382, 24'd7866452, 24'd8141855, 
24'd8466090, 24'd8774992, 24'd9007428, 24'd9117402, 24'd9083148, 24'd8911446, 24'd8636275, 24'd8312091, 24'd8003050, 24'd7770310, 24'd7659930, 24'd7693753, 24'd7865088, 24'd8140025, 24'd8464157, 24'd8773338, 24'd9006381, 24'd9117168, 24'd9083774, 24'd8912808, 24'd8638104, 24'd8314025, 24'd8004705, 24'd7771359, 24'd7660166, 24'd7693130, 24'd7863727, 24'd8138197, 24'd8462224, 24'd8771681, 
24'd9005329, 24'd9116929, 24'd9084395, 24'd8914167, 24'd8639931, 24'd8315958, 24'd8006363, 24'd7772413, 24'd7660407, 24'd7692511, 24'd7862370, 24'd8136371, 24'd8460290, 24'd8770022, 24'd9004273, 24'd9116685, 24'd9085012, 24'd8915522, 24'd8641756, 24'd8317893, 24'd8008024, 24'd7773472, 24'd7660654, 24'd7691897, 24'd7861017, 24'd8134547, 24'd8458355, 24'd8768360, 24'd9003213, 24'd9116436, 
24'd9085624, 24'd8916873, 24'd8643579, 24'd8319827, 24'd8009687, 24'd7774534, 24'd7660905, 24'd7691287, 24'd7859668, 24'd8132725, 24'd8456420, 24'd8766695, 24'd9002148, 24'd9116182, 24'd9086230, 24'd8918220, 24'd8645401, 24'd8321763, 24'd8011353, 24'd7775601, 24'd7661162, 24'd7690683, 24'd7858322, 24'd8130904, 24'd8454484, 24'd8765028, 24'd9001079, 24'd9115923, 24'd9086832, 24'd8919564, 
24'd8647221, 24'd8323698, 24'd8013021, 24'd7776672, 24'd7661424, 24'd7690084, 24'd7856980, 24'd8129085, 24'd8452548, 24'd8763358, 24'd9000006, 24'd9115658, 24'd9087429, 24'd8920904, 24'd8649039, 24'd8325635, 24'd8014693, 24'd7777748, 24'd7661691, 24'd7689489, 24'd7855642, 24'd8127268, 24'd8450612, 24'd8761686, 24'd8998928, 24'd9115389, 24'd9088021, 24'd8922241, 24'd8650855, 24'd8327571, 
24'd8016366, 24'd7778827, 24'd7661963, 24'd7688900, 24'd7854307, 24'd8125452, 24'd8448675, 24'd8760011, 24'd8997846, 24'd9115115, 24'd9088608, 24'd8923573, 24'd8652670, 24'd8329508, 24'd8018043, 24'd7779911, 24'd7662240, 24'd7688315, 24'd7852977, 24'd8123639, 24'd8446738, 24'd8758333, 24'd8996760, 24'd9114835, 24'd9089191, 24'd8924902, 24'd8654482, 24'd8331446, 24'd8019722, 24'd7781000, 
24'd7662522, 24'd7687735, 24'd7851650, 24'd8121827, 24'd8444800, 24'd8756653, 24'd8995670, 24'd9114550, 24'd9089768, 24'd8926227, 24'd8656293, 24'd8333384, 24'd8021403, 24'd7782092, 24'd7662809, 24'd7687160, 24'd7850327, 24'd8120018, 24'd8442862, 24'd8754970, 24'd8994575, 24'd9114260, 24'd9090340, 24'd8927549, 24'd8658102, 24'd8335322, 24'd8023088, 24'd7783189, 24'd7663101, 24'd7686590, 
24'd7849007, 24'd8118210, 24'd8440924, 24'd8753284, 24'd8993476, 24'd9113966, 24'd9090908, 24'd8928866, 24'd8659908, 24'd8337261, 24'd8024774, 24'd7784290, 24'd7663399, 24'd7686025, 24'd7847691, 24'd8116404, 24'd8438985, 24'd8751596, 24'd8992373, 24'd9113666, 24'd9091470, 24'd8930180, 24'd8661713, 24'd8339200, 24'd8026464, 24'd7785395, 24'd7663701, 24'd7685465, 24'd7846380, 24'd8114600, 
24'd8437046, 24'd8749906, 24'd8991266, 24'd9113361, 24'd9092028, 24'd8931490, 24'd8663516, 24'd8341139, 24'd8028155, 24'd7786505, 24'd7664009, 24'd7684910, 24'd7845071, 24'd8112798, 24'd8435106, 24'd8748213, 24'd8990154, 24'd9113050, 24'd9092581, 24'd8932796, 24'd8665318, 24'd8343079, 24'd8029850, 24'd7787618, 24'd7664322, 24'd7684360, 24'd7843767, 24'd8110998, 24'd8433166, 24'd8746517, 
24'd8989038, 24'd9112735, 24'd9093129, 24'd8934099, 24'd8667117, 24'd8345019, 24'd8031547, 24'd7788736, 24'd7664639, 24'd7683814, 24'd7842467, 24'd8109199, 24'd8431226, 24'd8744819, 24'd8987918, 24'd9112415, 24'd9093671, 24'd8935397, 24'd8668914, 24'd8346959, 24'd8033246, 24'd7789858, 24'd7664962, 24'd7683274, 24'd7841170, 24'd8107403, 24'd8429286, 24'd8743118, 24'd8986794, 24'd9112090, 
24'd9094209, 24'd8936692, 24'd8670709, 24'd8348899, 24'd8034948, 24'd7790985, 24'd7665290, 24'd7682739, 24'd7839877, 24'd8105609, 24'd8427345, 24'd8741415, 24'd8985666, 24'd9111759, 24'd9094742, 24'd8937983, 24'd8672503, 24'd8350840, 24'd8036652, 24'd7792115, 24'd7665623, 24'd7682208, 24'd7838588, 24'd8103816, 24'd8425404, 24'd8739710, 24'd8984533, 24'd9111424, 24'd9095270, 24'd8939270, 
24'd8674294, 24'd8352781, 24'd8038359, 24'd7793250, 24'd7665961, 24'd7681683, 24'd7837303, 24'd8102026, 24'd8423463, 24'd8738002, 24'd8983396, 24'd9111083, 24'd9095793, 24'd8940553, 24'd8676083, 24'd8354723, 24'd8040068, 24'd7794389, 24'd7666304, 24'd7681162, 24'd7836022, 24'd8100238, 24'd8421521, 24'd8736291, 24'd8982255, 24'd9110737, 24'd9096311, 24'd8941832, 24'd8677871, 24'd8356664, 
24'd8041780, 24'd7795532, 24'd7666652, 24'd7680646, 24'd7834745, 24'd8098452, 24'd8419580, 24'd8734578, 24'd8981110, 24'd9110387, 24'd9096825, 24'd8943107, 24'd8679656, 24'd8358606, 24'd8043494, 24'd7796679, 24'd7667006, 24'd7680136, 24'd7833471, 24'd8096667, 24'd8417638, 24'd8732863, 24'd8979961, 24'd9110031, 24'd9097333, 24'd8944379, 24'd8681439, 24'd8360548, 24'd8045211, 24'd7797830, 
24'd7667364, 24'd7679630, 24'd7832202, 24'd8094885, 24'd8415696, 24'd8731145, 24'd8978807, 24'd9109670, 24'd9097836, 24'd8945647, 24'd8683220, 24'd8362491, 24'd8046929, 24'd7798986, 24'd7667727, 24'd7679129, 24'd7830936, 24'd8093105, 24'd8413753, 24'd8729425, 24'd8977650, 24'd9109304, 24'd9098334, 24'd8946910, 24'd8684999, 24'd8364433, 24'd8048651, 24'd7800145, 24'd7668096, 24'd7678634, 
24'd7829674, 24'd8091327, 24'd8411811, 24'd8727703, 24'd8976488, 24'd9108933, 24'd9098827, 24'd8948170, 24'd8686776, 24'd8366376, 24'd8050375, 24'd7801309, 24'd7668469, 24'd7678143, 24'd7828417, 24'd8089551, 24'd8409868, 24'd8725978, 24'd8975322, 24'd9108557, 24'd9099316, 24'd8949426, 24'd8688551, 24'd8368318, 24'd8052101, 24'd7802477, 24'd7668848, 24'd7677657, 24'd7827163, 24'd8087777, 
24'd8407925, 24'd8724250, 24'd8974152, 24'd9108176, 24'd9099799, 24'd8950678, 24'd8690324, 24'd8370261, 24'd8053829, 24'd7803649, 24'd7669231, 24'd7677176, 24'd7825913, 24'd8086005, 24'd8405982, 24'd8722521, 24'd8972978, 24'd9107790, 24'd9100277, 24'd8951926, 24'd8692095, 24'd8372204, 24'd8055560, 24'd7804825, 24'd7669620, 24'd7676701, 24'd7824667, 24'd8084236, 24'd8404039, 24'd8720789, 
24'd8971800, 24'd9107399, 24'd9100750, 24'd8953170, 24'd8693864, 24'd8374148, 24'd8057293, 24'd7806005, 24'd7670013, 24'd7676230, 24'd7823425, 24'd8082468, 24'd8402096, 24'd8719054, 24'd8970618, 24'd9107003, 24'd9101219, 24'd8954410, 24'd8695630, 24'd8376091, 24'd8059029, 24'd7807190, 24'd7670412, 24'd7675764, 24'd7822186, 24'd8080703, 24'd8400153, 24'd8717318, 24'd8969432, 24'd9106602, 
24'd9101682, 24'd8955646, 24'd8697394, 24'd8378034, 24'd8060766, 24'd7808378, 24'd7670816, 24'd7675303, 24'd7820952, 24'd8078939, 24'd8398209, 24'd8715579, 24'd8968241, 24'd9106196, 24'd9102140, 24'd8956878, 24'd8699156, 24'd8379978, 24'd8062506, 24'd7809570, 24'd7671224, 24'd7674847, 24'd7819722, 24'd8077178, 24'd8396266, 24'd8713838, 24'd8967047, 24'd9105784, 24'd9102594, 24'd8958106, 
24'd8700916, 24'd8381921, 24'd8064249, 24'd7810767, 24'd7671638, 24'd7674397, 24'd7818496, 24'd8075419, 24'd8394322, 24'd8712094, 24'd8965849, 24'd9105368, 24'd9103042, 24'd8959331, 24'd8702674, 24'd8383865, 24'd8065994, 24'd7811967, 24'd7672057, 24'd7673951, 24'd7817274, 24'd8073663, 24'd8392379, 24'd8710348, 24'd8964646, 24'd9104947, 24'd9103485, 24'd8960551, 24'd8704430, 24'd8385808, 
24'd8067740, 24'd7813172, 24'd7672481, 24'd7673510, 24'd7816056, 24'd8071908, 24'd8390435, 24'd8708600, 24'd8963439, 24'd9104520, 24'd9103924, 24'd8961767, 24'd8706183, 24'd8387752, 24'd8069490, 24'd7814380, 24'd7672910, 24'd7673074, 24'd7814842, 24'd8070156, 24'd8388492, 24'd8706850, 24'd8962229, 24'd9104089, 24'd9104357, 24'd8962979, 24'd8707934, 24'd8389695, 24'd8071241, 24'd7815593, 
24'd7673344, 24'd7672643, 24'd7813631, 24'd8068406, 24'd8386548, 24'd8705097, 24'd8961014, 24'd9103653, 24'd9104785, 24'd8964187, 24'd8709683, 24'd8391639, 24'd8072995, 24'd7816810, 24'd7673782, 24'd7672218, 24'd7812425, 24'd8066658, 24'd8384604, 24'd8703343, 24'd8959796, 24'd9103211, 24'd9105208, 24'd8965391, 24'd8711430, 24'd8393582, 24'd8074750, 24'd7818030, 24'd7674226, 24'd7671797, 
24'd7811223, 24'd8064913, 24'd8382661, 24'd8701586, 24'd8958573, 24'd9102765, 24'd9105626, 24'd8966591, 24'd8713174, 24'd8395526, 24'd8076508, 24'd7819255, 24'd7674675, 24'd7671381, 24'd7810025, 24'd8063170, 24'd8380717, 24'd8699827, 24'd8957346, 24'd9102314, 24'd9106040, 24'd8967787, 24'd8714916, 24'd8397469, 24'd8078269, 24'd7820484, 24'd7675129, 24'd7670971, 24'd7808831, 24'd8061429, 
24'd8378774, 24'd8698065, 24'd8956116, 24'd9101857, 24'd9106448, 24'd8968979, 24'd8716656, 24'd8399413, 24'd8080031, 24'd7821716, 24'd7675588, 24'd7670565, 24'd7807641, 24'd8059690, 24'd8376831, 24'd8696302, 24'd8954881, 24'd9101396, 24'd9106851, 24'd8970167, 24'd8718394, 24'd8401356, 24'd8081796, 24'd7822953, 24'd7676052, 24'd7670164, 24'd7806456, 24'd8057954, 24'd8374887, 24'd8694536, 
24'd8953642, 24'd9100929, 24'd9107249, 24'd8971351, 24'd8720129, 24'd8403299, 24'd8083562, 24'd7824193, 24'd7676521, 24'd7669769, 24'd7805274, 24'd8056220, 24'd8372944, 24'd8692768, 24'd8952400, 24'd9100458, 24'd9107642, 24'd8972530, 24'd8721862, 24'd8405242, 24'd8085331, 24'd7825438, 24'd7676995, 24'd7669378, 24'd7804096, 24'd8054488, 24'd8371001, 24'd8690999, 24'd8951153, 24'd9099982, 
24'd9108030, 24'd8973706, 24'd8723592, 24'd8407185, 24'd8087102, 24'd7826686, 24'd7677474, 24'd7668993, 24'd7802923, 24'd8052758, 24'd8369058, 24'd8689227, 24'd8949903, 24'd9099500, 24'd9108413, 24'd8974877, 24'd8725320, 24'd8409128, 24'd8088875, 24'd7827939, 24'd7677957, 24'd7668613, 24'd7801753, 24'd8051031, 24'd8367115, 24'd8687452, 24'd8948649, 24'd9099014, 24'd9108791, 24'd8976045, 
24'd8727046, 24'd8411071, 24'd8090650, 24'd7829195, 24'd7678446, 24'd7668237, 24'd7800588, 24'd8049307, 24'd8365173, 24'd8685676, 24'd8947390, 24'd9098522, 24'd9109164, 24'd8977208, 24'd8728770, 24'd8413014, 24'd8092428, 24'd7830455, 24'd7678940, 24'd7667867, 24'd7799427, 24'd8047585, 24'd8363230, 24'd8683898, 24'd8946128, 24'd9098026, 24'd9109531, 24'd8978367, 24'd8730491, 24'd8414956, 
24'd8094207, 24'd7831719, 24'd7679439, 24'd7667502, 24'd7798270, 24'd8045865, 24'd8361288, 24'd8682117, 24'd8944862, 24'd9097525, 24'd9109894, 24'd8979522, 24'd8732209, 24'd8416898, 24'd8095989, 24'd7832988, 24'd7679943, 24'd7667141, 24'd7797117, 24'd8044147, 24'd8359346, 24'd8680335, 24'd8943592, 24'd9097019, 24'd9110252, 24'd8980673, 24'd8733926, 24'd8418840, 24'd8097772, 24'd7834259, 
24'd7680451, 24'd7666786, 24'd7795968, 24'd8042432, 24'd8357404, 24'd8678550, 24'd8942318, 24'd9096507, 24'd9110605, 24'd8981820, 24'd8735639, 24'd8420782, 24'd8099558, 24'd7835535, 24'd7680965, 24'd7666436, 24'd7794823, 24'd8040720, 24'd8355462, 24'd8676764, 24'd8941040, 24'd9095991, 24'd9110952, 24'd8982962, 24'd8737351, 24'd8422724, 24'd8101345, 24'd7836815, 24'd7681484, 24'd7666091, 
24'd7793683, 24'd8039009, 24'd8353521, 24'd8674975, 24'd8939759, 24'd9095470, 24'd9111295, 24'd8984101, 24'd8739060, 24'd8424665, 24'd8103135, 24'd7838099, 24'd7682007, 24'd7665751, 24'd7792547, 24'd8037302, 24'd8351579, 24'd8673185, 24'd8938473, 24'd9094944, 24'd9111632, 24'd8985235, 24'd8740766, 24'd8426606, 24'd8104926, 24'd7839386, 24'd7682536, 24'd7665416, 24'd7791415, 24'd8035596, 
24'd8349638, 24'd8671392, 24'd8937184, 24'd9094413, 24'd9111964, 24'd8986365, 24'd8742470, 24'd8428547, 24'd8106720, 24'd7840677, 24'd7683070, 24'd7665086, 24'd7790287, 24'd8033894, 24'd8347698, 24'd8669598, 24'd8935890, 24'd9093877, 24'd9112292, 24'd8987491, 24'd8744172, 24'd8430488, 24'd8108515, 24'd7841973, 24'd7683608, 24'd7664762, 24'd7789163, 24'd8032193, 24'd8345757, 24'd8667801, 
24'd8934593, 24'd9093336, 24'd9112614, 24'd8988612, 24'd8745871, 24'd8432428, 24'd8110313, 24'd7843272, 24'd7684151, 24'd7664442, 24'd7788043, 24'd8030495, 24'd8343817, 24'd8666003, 24'd8933292, 24'd9092790, 24'd9112931, 24'd8989730, 24'd8747568, 24'd8434368, 24'd8112112, 24'd7844574, 24'd7684700, 24'd7664127, 24'd7786928, 24'd8028800, 24'd8341877, 24'd8664202, 24'd8931988, 24'd9092239, 
24'd9113243, 24'd8990843, 24'd8749262, 24'd8436307, 24'd8113914, 24'd7845881, 24'd7685253, 24'd7663818, 24'd7785817, 24'd8027107, 24'd8339938, 24'd8662400, 24'd8930679, 24'd9091683, 24'd9113550, 24'd8991952, 24'd8750953, 24'd8438247, 24'd8115717, 24'd7847192, 24'd7685811, 24'd7663513, 24'd7784710, 24'd8025417, 24'd8337999, 24'd8660596, 24'd8929367, 24'd9091123, 24'd9113852, 24'd8993057, 
24'd8752642, 24'd8440186, 24'd8117522, 24'd7848506, 24'd7686375, 24'd7663214, 24'd7783607, 24'd8023729, 24'd8336060, 24'd8658790, 24'd8928051, 24'd9090557, 24'd9114149, 24'd8994157, 24'd8754329, 24'd8442124, 24'd8119329, 24'd7849824, 24'd7686943, 24'd7662920, 24'd7782509, 24'd8022044, 24'd8334122, 24'd8656982, 24'd8926731, 24'd9089986, 24'd9114441, 24'd8995254, 24'd8756012, 24'd8444063, 
24'd8121138, 24'd7851146, 24'd7687516, 24'd7662631, 24'd7781415, 24'd8020362, 24'd8332184, 24'd8655172, 24'd8925407, 24'd9089411, 24'd9114727, 24'd8996346, 24'd8757694, 24'd8446000, 24'd8122949, 24'd7852471, 24'd7688094, 24'd7662346, 24'd7780325, 24'd8018682, 24'd8330246, 24'd8653360, 24'd8924080, 24'd9088831, 24'd9115009, 24'd8997433, 24'd8759372, 24'd8447938, 24'd8124762, 24'd7853800, 
24'd7688676, 24'd7662067, 24'd7779239, 24'd8017004, 24'd8328309, 24'd8651546, 24'd8922749, 24'd9088245, 24'd9115285, 24'd8998517, 24'd8761048, 24'd8449875, 24'd8126576, 24'd7855134, 24'd7689264, 24'd7661794, 24'd7778158, 24'd8015329, 24'd8326372, 24'd8649731, 24'd8921414, 24'd9087655, 24'd9115556, 24'd8999596, 24'd8762722, 24'd8451811, 24'd8128393, 24'd7856470, 24'd7689857, 24'd7661525, 
24'd7777081, 24'd8013657, 24'd8324436, 24'd8647913, 24'd8920075, 24'd9087060, 24'd9115823, 24'd9000671, 24'd8764393, 24'd8453747, 24'd8130211, 24'd7857811, 24'd7690454, 24'd7661261, 24'd7776008, 24'd8011988, 24'd8322500, 24'd8646094, 24'd8918732, 24'd9086460, 24'd9116084, 24'd9001742, 24'd8766061, 24'd8455683, 24'd8132031, 24'd7859155, 24'd7691057, 24'd7661002, 24'd7774940, 24'd8010321, 
24'd8320564, 24'd8644273, 24'd8917386, 24'd9085855, 24'd9116340, 24'd9002808, 24'd8767727, 24'd8457618, 24'd8133853, 24'd7860503, 24'd7691664, 24'd7660749, 24'd7773876, 24'd8008657, 24'd8318629, 24'd8642450, 24'd8916037, 24'd9085245, 24'd9116591, 24'd9003870, 24'd8769390, 24'd8459553, 24'd8135677, 24'd7861855, 24'd7692276, 24'd7660500, 24'd7772816, 24'd8006995, 24'd8316695, 24'd8640626, 
24'd8914683, 24'd9084631, 24'd9116837, 24'd9004928, 24'd8771050, 24'd8461487, 24'd8137502, 24'd7863210, 24'd7692893, 24'd7660257, 24'd7771760, 24'd8005336, 24'd8314761, 24'd8638800, 24'd8913326, 24'd9084011, 24'd9117078, 24'd9005981, 24'd8772707, 24'd8463421, 24'd8139329, 24'd7864569, 24'd7693515, 24'd7660019, 24'd7770709, 24'd8003680, 24'd8312827, 24'd8636971, 24'd8911965, 24'd9083387, 
24'd9117313, 24'd9007030, 24'd8774362, 24'd8465354, 24'd8141158, 24'd7865932, 24'd7694142, 24'd7659786, 24'd7769662, 24'd8002026, 24'd8310894, 24'd8635142, 24'd8910600, 24'd9082758, 24'd9117544, 24'd9008075, 24'd8776014, 24'd8467287, 24'd8142989, 24'd7867298, 24'd7694774, 24'd7659558, 24'd7768619, 24'd8000376, 24'd8308962, 24'd8633310, 24'd8909232, 24'd9082123, 24'd9117769, 24'd9009115, 
24'd8777664, 24'd8469219, 24'd8144821, 24'd7868668, 24'd7695411, 24'd7659335, 24'd7767581, 24'd7998727, 24'd8307030, 24'd8631477, 24'd8907860, 24'd9081484, 24'd9117989, 24'd9010151, 24'd8779311, 24'd8471151, 24'd8146655, 24'd7870042, 24'd7696052, 24'd7659117, 24'd7766547, 24'd7997082, 24'd8305099, 24'd8629642, 24'd8906485, 24'd9080840, 24'd9118205, 24'd9011183, 24'd8780955, 24'd8473081, 
24'd8148491, 24'd7871419, 24'd7696698, 24'd7658905, 24'd7765518, 24'd7995439, 24'd8303168, 24'd8627805, 24'd8905106, 24'd9080192, 24'd9118415, 24'd9012210, 24'd8782596, 24'd8475012, 24'd8150329, 24'd7872800, 24'd7697349, 24'd7658697, 24'd7764493, 24'd7993800, 24'd8301238, 24'd8625967, 24'd8903723, 24'd9079538, 24'd9118620, 24'd9013233, 24'd8784234, 24'd8476942, 24'd8152168, 24'd7874185, 
24'd7698005, 24'd7658495, 24'd7763472, 24'd7992163, 24'd8299309, 24'd8624127, 24'd8902336, 24'd9078880, 24'd9118820, 24'd9014252, 24'd8785870, 24'd8478871, 24'd8154009, 24'd7875573, 24'd7698666, 24'd7658297, 24'd7762456, 24'd7990528, 24'd8297380, 24'd8622285, 24'd8900946, 24'd9078217, 24'd9119014, 24'd9015266, 24'd8787503, 24'd8480799, 24'd8155851, 24'd7876965, 24'd7699332, 24'd7658105, 
24'd7761444, 24'd7988897, 24'd8295452, 24'd8620442, 24'd8899553, 24'd9077548, 24'd9119204, 24'd9016276, 24'd8789133, 24'd8482727, 24'd8157695, 24'd7878360, 24'd7700002, 24'd7657918, 24'd7760436, 24'd7987268, 24'd8293524, 24'd8618597, 24'd8898156, 24'd9076876, 24'd9119388, 24'd9017281, 24'd8790760, 24'd8484654, 24'd8159541, 24'd7879759, 24'd7700678, 24'd7657736, 24'd7759433, 24'd7985642, 
24'd8291597, 24'd8616751, 24'd8896755, 24'd9076198, 24'd9119568, 24'd9018282, 24'd8792385, 24'd8486581, 24'd8161388, 24'd7881162, 24'd7701358, 24'd7657560, 24'd7758434, 24'd7984019, 24'd8289671, 24'd8614903, 24'd8895351, 24'd9075515, 24'd9119742, 24'd9019279, 24'd8794006, 24'd8488507, 24'd8163237, 24'd7882568, 24'd7702043, 24'd7657388, 24'd7757440, 24'd7982399, 24'd8287746, 24'd8613053, 
24'd8893943, 24'd9074828, 24'd9119911, 24'd9020271, 24'd8795625, 24'd8490432, 24'd8165088, 24'd7883977, 24'd7702733, 24'd7657221, 24'd7756450, 24'd7980781, 24'd8285821, 24'd8611202, 24'd8892531, 24'd9074136, 24'd9120075, 24'd9021258, 24'd8797241, 24'd8492356, 24'd8166940, 24'd7885391, 24'd7703427, 24'd7657060, 24'd7755464, 24'd7979167, 24'd8283897, 24'd8609349, 24'd8891117, 24'd9073439, 
24'd9120234, 24'd9022242, 24'd8798854, 24'd8494280, 24'd8168793, 24'd7886807, 24'd7704127, 24'd7656904, 24'd7754483, 24'd7977555, 24'd8281973, 24'd8607494, 24'd8889698, 24'd9072737, 24'd9120388, 24'd9023220, 24'd8800465, 24'd8496203, 24'd8170648, 24'd7888227, 24'd7704831, 24'd7656752, 24'd7753507, 24'd7975946, 24'd8280051, 24'd8605639, 24'd8888276, 24'd9072030, 24'd9120536, 24'd9024195, 
24'd8802072, 24'd8498125, 24'd8172505, 24'd7889651, 24'd7705540, 24'd7656606, 24'd7752535, 24'd7974341, 24'd8278129, 24'd8603781, 24'd8886851, 24'd9071319, 24'd9120680, 24'd9025165, 24'd8803676, 24'd8500047, 24'd8174363, 24'd7891078, 24'd7706254, 24'd7656466, 24'd7751567, 24'd7972738, 24'd8276208, 24'd8601922, 24'd8885422, 24'd9070603, 24'd9120818, 24'd9026130, 24'd8805278, 24'd8501967, 
24'd8176223, 24'd7892509, 24'd7706972, 24'd7656330, 24'd7750604, 24'd7971138, 24'd8274288, 24'd8600062, 24'd8883989, 24'd9069882, 24'd9120951, 24'd9027091, 24'd8806876, 24'd8503887, 24'd8178084, 24'd7893943, 24'd7707696, 24'd7656199, 24'd7749645, 24'd7969540, 24'd8272368, 24'd8598200, 24'd8882553, 24'd9069156, 24'd9121079, 24'd9028048, 24'd8808472, 24'd8505806, 24'd8179947, 24'd7895381, 
24'd7708424, 24'd7656074, 24'd7748691, 24'd7967946, 24'd8270450, 24'd8596336, 24'd8881114, 24'd9068425, 24'd9121202, 24'd9029000, 24'd8810065, 24'd8507724, 24'd8181811, 24'd7896822, 24'd7709157, 24'd7655953, 24'd7747741, 24'd7966355, 24'd8268532, 24'd8594472, 24'd8879671, 24'd9067690, 24'd9121320, 24'd9029947, 24'd8811655, 24'd8509642, 24'd8183676, 24'd7898267, 24'd7709894, 24'd7655838, 
24'd7746796, 24'd7964767, 24'd8266615, 24'd8592605, 24'd8878225, 24'd9066950, 24'd9121433, 24'd9030890, 24'd8813241, 24'd8511558, 24'd8185543, 24'd7899715, 24'd7710637, 24'd7655728, 24'd7745855, 24'd7963181, 24'd8264699, 24'd8590738, 24'd8876775, 24'd9066205, 24'd9121540, 24'd9031829, 24'd8814825, 24'd8513474, 24'd8187412, 24'd7901166, 24'd7711384, 24'd7655623, 24'd7744919, 24'd7961599, 
24'd8262784, 24'd8588868, 24'd8875322, 24'd9065456, 24'd9121642, 24'd9032763, 24'd8816406, 24'd8515389, 24'd8189282, 24'd7902621, 24'd7712136, 24'd7655523, 24'd7743987, 24'd7960020, 24'd8260869, 24'd8586998, 24'd8873866, 24'd9064701, 24'd9121740, 24'd9033692, 24'd8817984, 24'd8517303, 24'd8191153, 24'd7904079, 24'd7712892, 24'd7655429, 24'd7743060, 24'd7958443, 24'd8258956, 24'd8585126, 
24'd8872406, 24'd9063942, 24'd9121832, 24'd9034617, 24'd8819559, 24'd8519216, 24'd8193026, 24'd7905541, 24'd7713654, 24'd7655339, 24'd7742137, 24'd7956870, 24'd8257043, 24'd8583253, 24'd8870942, 24'd9063179, 24'd9121919, 24'd9035538, 24'd8821131, 24'd8521128, 24'd8194900, 24'd7907006, 24'd7714420, 24'd7655255, 24'd7741219, 24'd7955300, 24'd8255132, 24'd8581378, 24'd8869476, 24'd9062410, 
24'd9122000, 24'd9036454, 24'd8822699, 24'd8523039, 24'd8196775, 24'd7908474, 24'd7715191, 24'd7655176, 24'd7740305, 24'd7953732, 24'd8253221, 24'd8579502, 24'd8868005, 24'd9061637, 24'd9122077, 24'd9037365, 24'd8824265, 24'd8524949, 24'd8198652, 24'd7909946, 24'd7715966, 24'd7655101, 24'd7739396, 24'd7952168, 24'd8251311, 24'd8577625, 24'd8866532, 24'd9060859, 24'd9122149, 24'd9038272, 
24'd8825828, 24'd8526858, 24'd8200530, 24'd7911421, 24'd7716747, 24'd7655032, 24'd7738491, 24'd7950607, 24'd8249402, 24'd8575746, 24'd8865055, 24'd9060076, 24'd9122215, 24'd9039174, 24'd8827387, 24'd8528767, 24'd8202409, 24'd7912899, 24'd7717532, 24'd7654969, 24'd7737591, 24'd7949049, 24'd8247494, 24'd8573866, 24'd8863575, 24'd9059289, 24'd9122276, 24'd9040072, 24'd8828944, 24'd8530674, 
24'd8204290, 24'd7914381, 24'd7718321, 24'd7654910, 24'd7736696, 24'd7947494, 24'd8245588, 24'd8571985, 24'd8862092, 24'd9058497, 24'd9122332, 24'd9040965, 24'd8830497, 24'd8532580, 24'd8206172, 24'd7915866, 24'd7719116, 24'd7654857, 24'd7735805, 24'd7945942, 24'd8243682, 24'd8570102, 24'd8860605, 24'd9057700, 24'd9122383, 24'd9041854, 24'd8832048, 24'd8534486, 24'd8208055, 24'd7917355, 
24'd7719915, 24'd7654808, 24'd7734919, 24'd7944393, 24'd8241777, 24'd8568218, 24'd8859115, 24'd9056899, 24'd9122429, 24'd9042738, 24'd8833595, 24'd8536390, 24'd8209939, 24'd7918847, 24'd7720719, 24'd7654765, 24'd7734037, 24'd7942848, 24'd8239873, 24'd8566333, 24'd8857621, 24'd9056093, 24'd9122470, 24'd9043617, 24'd8835139, 24'd8538293, 24'd8211825, 24'd7920342, 24'd7721527, 24'd7654727, 
24'd7733160, 24'd7941305, 24'd8237970, 24'd8564447, 24'd8856125, 24'd9055282, 24'd9122505, 24'd9044492, 24'd8836680, 24'd8540195, 24'd8213712, 24'd7921840, 24'd7722340, 24'd7654694, 24'd7732288, 24'd7939766, 24'd8236069, 24'd8562559, 24'd8854625, 24'd9054466, 24'd9122536, 24'd9045362, 24'd8838218, 24'd8542097, 24'd8215600, 24'd7923342, 24'd7723158, 24'd7654666, 24'd7731420, 24'd7938229, 
24'd8234168, 24'd8560670, 24'd8853121, 24'd9053646, 24'd9122561, 24'd9046228, 24'd8839753, 24'd8543997, 24'd8217490, 24'd7924846, 24'd7723981, 24'd7654643, 24'd7730556, 24'd7936696, 24'd8232269, 24'd8558780, 24'd8851615, 24'd9052821, 24'd9122581, 24'd9047089, 24'd8841284, 24'd8545896, 24'd8219380, 24'd7926355, 24'd7724808, 24'd7654626, 24'd7729698, 24'd7935166, 24'd8230370, 24'd8556889, 
24'd8850105, 24'd9051992, 24'd9122596, 24'd9047945, 24'd8842812, 24'd8547794, 24'd8221272, 24'd7927866, 24'd7725640, 24'd7654614, 24'd7728844, 24'd7933640, 24'd8228473, 24'd8554997, 24'd8848592, 24'd9051158, 24'd9122606, 24'd9048797, 24'd8844338, 24'd8549690, 24'd8223165, 24'd7929380, 24'd7726476, 24'd7654606, 24'd7727994, 24'd7932116, 24'd8226577, 24'd8553103, 24'd8847076, 24'd9050319, 
24'd9122610, 24'd9049644, 24'd8845860, 24'd8551586, 24'd8225059, 24'd7930898, 24'd7727317, 24'd7654604, 24'd7727149, 24'd7930596, 24'd8224682, 24'd8551208, 24'd8845557, 24'd9049475, 24'd9122610, 24'd9050486, 24'd8847378, 24'd8553480, 24'd8226954, 24'd7932419, 24'd7728163, 24'd7654607, 24'd7726309, 24'd7929078, 24'd8222788, 24'd8549312, 24'd8844034, 24'd9048627, 24'd9122604, 24'd9051324, 
24'd8848894, 24'd8555374, 24'd8228851, 24'd7933944, 24'd7729013, 24'd7654616, 24'd7725474, 24'd7927565, 24'd8220895, 24'd8547415, 24'd8842508, 24'd9047775, 24'd9122593, 24'd9052157, 24'd8850406, 24'd8557266, 24'd8230748, 24'd7935471, 24'd7729868, 24'd7654629, 24'd7724643, 24'd7926054, 24'd8219003, 24'd8545517, 24'd8840979, 24'd9046917, 24'd9122577, 24'd9052986, 24'd8851915, 24'd8559157, 
24'd8232647, 24'd7937002, 24'd7730728, 24'd7654648, 24'd7723816, 24'd7924546, 24'd8217113, 24'd8543618, 24'd8839447, 24'd9046056, 24'd9122556, 24'd9053810, 24'd8853421, 24'd8561047, 24'd8234547, 24'd7938535, 24'd7731592, 24'd7654671, 24'd7722995, 24'd7923042, 24'd8215224, 24'd8541718, 24'd8837912, 24'd9045189, 24'd9122530, 24'd9054629, 24'd8854924, 24'd8562935, 24'd8236448, 24'd7940072, 
24'd7732461, 24'd7654700, 24'd7722178, 24'd7921541, 24'd8213336, 24'd8539817, 24'd8836373, 24'd9044318, 24'd9122499, 24'd9055444, 24'd8856423, 24'd8564823, 24'd8238350, 24'd7941612, 24'd7733334, 24'd7654734, 24'd7721366, 24'd7920044, 24'd8211449, 24'd8537914, 24'd8834832, 24'd9043442, 24'd9122462, 24'd9056254, 24'd8857919, 24'd8566709, 24'd8240252, 24'd7943155, 24'd7734212, 24'd7654773, 
24'd7720558, 24'd7918549, 24'd8209564, 24'd8536011, 24'd8833287, 24'd9042562, 24'd9122420, 24'd9057059, 24'd8859412, 24'd8568594, 24'd8242156, 24'd7944702, 24'd7735095, 24'd7654817, 24'd7719755, 24'd7917058, 24'd8207679, 24'd8534106, 24'd8831739, 24'd9041677, 24'd9122374, 24'd9057859, 24'd8860901, 24'd8570477, 24'd8244061, 24'd7946251, 24'd7735982, 24'd7654867, 24'd7718957, 24'd7915570, 
24'd8205796, 24'd8532201, 24'd8830188, 24'd9040787, 24'd9122322, 24'd9058655, 24'd8862387, 24'd8572360, 24'd8245967, 24'd7947804, 24'd7736874, 24'd7654921, 24'd7718164, 24'd7914086, 24'd8203915, 24'd8530294, 24'd8828634, 24'd9039893, 24'd9122264, 24'd9059446, 24'd8863870, 24'd8574241, 24'd8247874, 24'd7949359, 24'd7737770, 24'd7654981, 24'd7717375, 24'd7912605, 24'd8202034, 24'd8528387, 
24'd8827077, 24'd9038995, 24'd9122202, 24'd9060233, 24'd8865350, 24'd8576120, 24'd8249783, 24'd7950918, 24'd7738671, 24'd7655046, 24'd7716591, 24'd7911127, 24'd8200155, 24'd8526478, 24'd8825517, 24'd9038092, 24'd9122135, 24'd9061014, 24'd8866826, 24'd8577999, 24'd8251691, 24'd7952480, 24'd7739577, 24'd7655116, 24'd7715812, 24'd7909652, 24'd8198278, 24'd8524569, 24'd8823953, 24'd9037184, 
24'd9122062, 24'd9061791, 24'd8868299, 24'd8579876, 24'd8253601, 24'd7954044, 24'd7740487, 24'd7655191, 24'd7715037, 24'd7908181, 24'd8196401, 24'd8522658, 24'd8822387, 24'd9036272, 24'd9121985, 24'd9062564, 24'd8869768, 24'd8581752, 24'd8255512, 24'd7955612, 24'd7741401, 24'd7655271, 24'd7714267, 24'd7906714, 24'd8194526, 24'd8520747, 24'd8820818, 24'd9035355, 24'd9121902, 24'd9063331, 
24'd8871234, 24'd8583626, 24'd8257424, 24'd7957183, 24'd7742320, 24'd7655357, 24'd7713502, 24'd7905249, 24'd8192652, 24'd8518835, 24'd8819245, 24'd9034433, 24'd9121814, 24'd9064094, 24'd8872697, 24'd8585499, 24'd8259337, 24'd7958757, 24'd7743244, 24'd7655447, 24'd7712741, 24'd7903788, 24'd8190780, 24'd8516921, 24'd8817670, 24'd9033507, 24'd9121721, 24'd9064852, 24'd8874156, 24'd8587371, 
24'd8261251, 24'd7960334, 24'd7744172, 24'd7655543, 24'd7711986, 24'd7902331, 24'd8188909, 24'd8515007, 24'd8816091, 24'd9032577, 24'd9121622, 24'd9065605, 24'd8875612, 24'd8589241, 24'd8263165, 24'd7961914, 24'd7745105, 24'd7655644, 24'd7711235, 24'd7900876, 24'd8187039, 24'd8513092, 24'd8814510, 24'd9031642, 24'd9121519, 24'd9066354, 24'd8877064, 24'd8591110, 24'd8265080, 24'd7963497, 
24'd7746042, 24'd7655750, 24'd7710488, 24'd7899426, 24'd8185171, 24'd8511176, 24'd8812925, 24'd9030703, 24'd9121411, 24'd9067098, 24'd8878513, 24'd8592977, 24'd8266997, 24'd7965083, 24'd7746984, 24'd7655861, 24'd7709747, 24'd7897978, 24'd8183305, 24'd8509260, 24'd8811338, 24'd9029759, 24'd9121297, 24'd9067837, 24'd8879959, 24'd8594843, 24'd8268914, 24'd7966672, 24'd7747930, 24'd7655977, 
24'd7709010, 24'd7896535, 24'd8181439, 24'd8507342, 24'd8809748, 24'd9028810, 24'd9121178, 24'd9068571, 24'd8881401, 24'd8596708, 24'd8270832, 24'd7968264, 24'd7748881, 24'd7656098, 24'd7708278, 24'd7895094, 24'd8179575, 24'd8505424, 24'd8808154, 24'd9027857, 24'd9121054, 24'd9069301, 24'd8882840, 24'd8598571, 24'd8272751, 24'd7969858, 24'd7749836, 24'd7656225, 24'd7707551, 24'd7893657, 
24'd8177713, 24'd8503505, 24'd8806558, 24'd9026900, 24'd9120925, 24'd9070026, 24'd8884275, 24'd8600433, 24'd8274670, 24'd7971456, 24'd7750795, 24'd7656356, 24'd7706829, 24'd7892224, 24'd8175852, 24'd8501585, 24'd8804959, 24'd9025938, 24'd9120791, 24'd9070746, 24'd8885707, 24'd8602293, 24'd8276591, 24'd7973057, 24'd7751759, 24'd7656493, 24'd7706111, 24'd7890794, 24'd8173993, 24'd8499664, 
24'd8803357, 24'd9024972, 24'd9120651, 24'd9071461, 24'd8887135, 24'd8604151, 24'd8278512, 24'd7974660, 24'd7752728, 24'd7656635, 24'd7705398, 24'd7889367, 24'd8172135, 24'd8497742, 24'd8801752, 24'd9024001, 24'd9120507, 24'd9072171, 24'd8888560, 24'd8606008, 24'd8280434, 24'd7976267, 24'd7753701, 24'd7656782, 24'd7704690, 24'd7887944, 24'd8170279, 24'd8495820, 24'd8800144, 24'd9023026, 
24'd9120357, 24'd9072877, 24'd8889981, 24'd8607864, 24'd8282357, 24'd7977876, 24'd7754679, 24'd7656934, 24'd7703987, 24'd7886525, 24'd8168424, 24'd8493897, 24'd8798533, 24'd9022046, 24'd9120203, 24'd9073578, 24'd8891399, 24'd8609718, 24'd8284280, 24'd7979488, 24'd7755660, 24'd7657092, 24'd7703289, 24'd7885109, 24'd8166570, 24'd8491973, 24'd8796919, 24'd9021062, 24'd9120043, 24'd9074274, 
24'd8892813, 24'd8611571, 24'd8286204, 24'd7981103, 24'd7756647, 24'd7657254, 24'd7702595, 24'd7883696, 24'd8164719, 24'd8490048, 24'd8795303, 24'd9020073, 24'd9119878, 24'd9074965, 24'd8894224, 24'd8613422, 24'd8288129, 24'd7982721, 24'd7757638, 24'd7657422, 24'd7701906, 24'd7882287, 24'd8162869, 24'd8488123, 24'd8793684, 24'd9019080, 24'd9119708, 24'd9075652, 24'd8895631, 24'd8615271, 
24'd8290055, 24'd7984342, 24'd7758633, 24'd7657594, 24'd7701222, 24'd7880882, 24'd8161020, 24'd8486197, 24'd8792061, 24'd9018083, 24'd9119532, 24'd9076333, 24'd8897034, 24'd8617119, 24'd8291981, 24'd7985966, 24'd7759633, 24'd7657772, 24'd7700543, 24'd7879480, 24'd8159173, 24'd8484270, 24'd8790436, 24'd9017081, 24'd9119352, 24'd9077010, 24'd8898434, 24'd8618965, 24'd8293908, 24'd7987592, 
24'd7760637, 24'd7657955, 24'd7699868, 24'd7878082, 24'd8157328, 24'd8482343, 24'd8788808, 24'd9016075, 24'd9119166, 24'd9077682, 24'd8899831, 24'd8620810, 24'd8295836, 24'd7989222, 24'd7761645, 24'd7658143, 24'd7699199, 24'd7876687, 24'd8155484, 24'd8480415, 24'd8787178, 24'd9015064, 24'd9118976, 24'd9078349, 24'd8901224, 24'd8622652, 24'd8297764, 24'd7990854, 24'd7762658, 24'd7658336, 
24'd7698534, 24'd7875296, 24'd8153642, 24'd8478486, 24'd8785544, 24'd9014049, 24'd9118780, 24'd9079011, 24'd8902613, 24'd8624494, 24'd8299693, 24'd7992489, 24'd7763675, 24'd7658535, 24'd7697874, 24'd7873909, 24'd8151801, 24'd8476557, 24'd8783908, 24'd9013030, 24'd9118579, 24'd9079669, 24'd8903999, 24'd8626333, 24'd8301623, 24'd7994126, 24'd7764697, 24'd7658738, 24'd7697219, 24'd7872525, 
24'd8149962, 24'd8474627, 24'd8782269, 24'd9012006, 24'd9118373, 24'd9080321, 24'd8905381, 24'd8628171, 24'd8303553, 24'd7995767, 24'd7765723, 24'd7658947, 24'd7696569, 24'd7871145, 24'd8148125, 24'd8472697, 24'd8780627, 24'd9010978, 24'd9118162, 24'd9080969, 24'd8906759, 24'd8630008, 24'd8305484, 24'd7997410, 24'd7766753, 24'd7659160, 24'd7695924, 24'd7869768, 24'd8146290, 24'd8470766, 
24'd8778983, 24'd9009945, 24'd9117946, 24'd9081612, 24'd8908134, 24'd8631842, 24'd8307415, 24'd7999056, 24'd7767788, 24'd7659379, 24'd7695283, 24'd7868395, 24'd8144456, 24'd8468834, 24'd8777335, 24'd9008908, 24'd9117725, 24'd9082250, 24'd8909505, 24'd8633675, 24'd8309347, 24'd8000704, 24'd7768827, 24'd7659603, 24'd7694648, 24'd7867026, 24'd8142624, 24'd8466902, 24'd8775685, 24'd9007867, 
24'd9117498, 24'd9082883, 24'd8910872, 24'd8635506, 24'd8311279, 24'd8002356, 24'd7769870, 24'd7659832, 24'd7694017, 24'd7865660, 24'd8140794, 24'd8464969, 24'd8774033, 24'd9006821, 24'd9117267, 24'd9083512, 24'd8912236, 24'd8637336, 24'd8313213, 24'd8004010, 24'd7770918, 24'd7660066, 24'd7693391, 24'd7864298, 24'd8138965, 24'd8463036, 24'd8772377, 24'd9005771, 24'd9117030, 24'd9084135, 
24'd8913596, 24'd8639164, 24'd8315146, 24'd8005666, 24'd7771970, 24'd7660305, 24'd7692770, 24'd7862940, 24'd8137138, 24'd8461102, 24'd8770719, 24'd9004717, 24'd9116788, 24'd9084754, 24'd8914953, 24'd8640990, 24'd8317080, 24'd8007326, 24'd7773027, 24'd7660550, 24'd7692154, 24'd7861585, 24'd8135313, 24'd8459168, 24'd8769058, 24'd9003659, 24'd9116541, 24'd9085367, 24'd8916306, 24'd8642814, 
24'd8319015, 24'd8008988, 24'd7774087, 24'd7660799, 24'd7691543, 24'd7860234, 24'd8133490, 24'd8457233, 24'd8767395, 24'd9002596, 24'd9116289, 24'd9085976, 24'd8917655, 24'd8644636, 24'd8320950, 24'd8010653, 24'd7775152, 24'd7661054, 24'd7690936, 24'd7858887, 24'd8131668, 24'd8455298, 24'd8765729, 24'd9001529, 24'd9116032, 24'd9086580, 24'd8919000, 24'd8646457, 24'd8322885, 24'd8012320, 
24'd7776222, 24'd7661313, 24'd7690335, 24'd7857543, 24'd8129849, 24'd8453362, 24'd8764060, 24'd9000457, 24'd9115770, 24'd9087179, 24'd8920342, 24'd8648276, 24'd8324821, 24'd8013990, 24'd7777295, 24'd7661578, 24'd7689738, 24'd7856204, 24'd8128031, 24'd8451426, 24'd8762389, 24'd8999381, 24'd9115503, 24'd9087773, 24'd8921680, 24'd8650093, 24'd8326758, 24'd8015663, 24'd7778373, 24'd7661848, 
24'd7689147, 24'd7854868, 24'd8126215, 24'd8449489, 24'd8760715, 24'd8998301, 24'd9115230, 24'd9088362, 24'd8923014, 24'd8651908, 24'd8328695, 24'd8017338, 24'd7779455, 24'd7662123, 24'd7688560, 24'd7853535, 24'd8124400, 24'd8447552, 24'd8759038, 24'd8997217, 24'd9114953, 24'd9088947, 24'd8924344, 24'd8653721, 24'd8330632, 24'd8019016, 24'd7780542, 24'd7662403, 24'd7687978, 24'd7852207, 
24'd8122588, 24'd8445614, 24'd8757359, 24'd8996128, 24'd9114670, 24'd9089526, 24'd8925671, 24'd8655532, 24'd8332570, 24'd8020697, 24'd7781633, 24'd7662688, 24'd7687401, 24'd7850882, 24'd8120778, 24'd8443676, 24'd8755677, 24'd8995035, 24'd9114383, 24'd9090101, 24'd8926994, 24'd8657342, 24'd8334508, 24'd8022380, 24'd7782728, 24'd7662978, 24'd7686829, 24'd7849561, 24'd8118969, 24'd8441738, 
24'd8753993, 24'd8993938, 24'd9114090, 24'd9090670, 24'd8928313, 24'd8659150, 24'd8336446, 24'd8024065, 24'd7783827, 24'd7663273, 24'd7686262, 24'd7848244, 24'd8117162, 24'd8439799, 24'd8752306, 24'd8992837, 24'd9113792, 24'd9091235, 24'd8929629, 24'd8660955, 24'd8338385, 24'd8025754, 24'd7784930, 24'd7663574, 24'd7685700, 24'd7846930, 24'd8115357, 24'd8437860, 24'd8750616, 24'd8991731, 
24'd9113489, 24'd9091794, 24'd8930940, 24'd8662759, 24'd8340324, 24'd8027444, 24'd7786038, 24'd7663879, 24'd7685143, 24'd7845620, 24'd8113554, 24'd8435921, 24'd8748924, 24'd8990622, 24'd9113181, 24'd9092349, 24'd8932248, 24'd8664561, 24'd8342264, 24'd8029138, 24'd7787150, 24'd7664190, 24'd7684590, 24'd7844315, 24'd8111753, 24'd8433981, 24'd8747230, 24'd8989507, 24'd9112868, 24'd9092899, 
24'd8933552, 24'd8666361, 24'd8344204, 24'd8030833, 24'd7788266, 24'd7664505, 24'd7684043, 24'd7843013, 24'd8109954, 24'd8432041, 24'd8745533, 24'd8988389, 24'd9112550, 24'd9093444, 24'd8934852, 24'd8668159, 24'd8346144, 24'd8032532, 24'd7789386, 24'd7664826, 24'd7683500, 24'd7841714, 24'd8108157, 24'd8430101, 24'd8743833, 24'd8987267, 24'd9112227, 24'd9093984, 24'd8936148, 24'd8669955, 
24'd8348084, 24'd8034233, 24'd7790511, 24'd7665152, 24'd7682963, 24'd7840420, 24'd8106362, 24'd8428160, 24'd8742131, 24'd8986140, 24'd9111899, 24'd9094519, 24'd8937441, 24'd8671750, 24'd8350025, 24'd8035936, 24'd7791640, 24'd7665483, 24'd7682430, 24'd7839129, 24'd8104569, 24'd8426219, 24'd8740427, 24'd8985009, 24'd9111565, 24'd9095049, 24'd8938729, 24'd8673542, 24'd8351966, 24'd8037642, 
24'd7792773, 24'd7665818, 24'd7681903, 24'd7837843, 24'd8102778, 24'd8424278, 24'd8738720, 24'd8983874, 24'd9111227, 24'd9095574, 24'd8940014, 24'd8675332, 24'd8353907, 24'd8039350, 24'd7793910, 24'd7666159, 24'd7681380, 24'd7836560, 24'd8100989, 24'd8422337, 24'd8737010, 24'd8982735, 24'd9110883, 24'd9096094, 24'd8941295, 24'd8677120, 24'd8355849, 24'd8041061, 24'd7795051, 24'd7666505, 
24'd7680862, 24'd7835281, 24'd8099202, 24'd8420395, 24'd8735298, 24'd8981592, 24'd9110535, 24'd9096610, 24'd8942572, 24'd8678906, 24'd8357791, 24'd8042774, 24'd7796197, 24'd7666857, 24'd7680350, 24'd7834006, 24'd8097416, 24'd8418453, 24'd8733584, 24'd8980444, 24'd9110181, 24'd9097120, 24'd8943845, 24'd8680690, 24'd8359733, 24'd8044489, 24'd7797346, 24'd7667213, 24'd7679842, 24'd7832735, 
24'd8095633, 24'd8416511, 24'd8731867, 24'd8979292, 24'd9109822, 24'd9097625, 24'd8945115, 24'd8682472, 24'd8361675, 24'd8046207, 24'd7798500, 24'd7667574, 24'd7679339, 24'd7831467, 24'd8093852, 24'd8414569, 24'd8730148, 24'd8978137, 24'd9109459, 24'd9098125, 24'd8946380, 24'd8684252, 24'd8363617, 24'd8047928, 24'd7799658, 24'd7667940, 24'd7678841, 24'd7830204, 24'd8092073, 24'd8412627, 
24'd8728426, 24'd8976977, 24'd9109090, 24'd9098621, 24'd8947641, 24'd8686030, 24'd8365560, 24'd8049650, 24'd7800820, 24'd7668312, 24'd7678348, 24'd7828944, 24'd8090297, 24'd8410684, 24'd8726702, 24'd8975813, 24'd9108716, 24'd9099111, 24'd8948899, 24'd8687806, 24'd8367502, 24'd8051375, 24'd7801986, 24'd7668688, 24'd7677861, 24'd7827689, 24'd8088522, 24'd8408741, 24'd8724976, 24'd8974644, 
24'd9108337, 24'd9099596, 24'd8950152, 24'd8689580, 24'd8369445, 24'd8053103, 24'd7803156, 24'd7669069, 24'd7677378, 24'd7826437, 24'd8086749, 24'd8406798, 24'd8723248, 24'd8973472, 24'd9107953, 24'd9100077, 24'd8951402, 24'd8691351, 24'd8371388, 24'd8054833, 24'd7804331, 24'd7669456, 24'd7676900, 24'd7825190, 24'd8084979, 24'd8404855, 24'd8721517, 24'd8972296, 24'd9107564, 24'd9100552, 
24'd8952648, 24'd8693121, 24'd8373331, 24'd8056565, 24'd7805509, 24'd7669847, 24'd7676427, 24'd7823946, 24'd8083210, 24'd8402912, 24'd8719783, 24'd8971115, 24'd9107170, 24'd9101023, 24'd8953890, 24'd8694888, 24'd8375275, 24'd8058299, 24'd7806692, 24'd7670244, 24'd7675959, 24'd7822706, 24'd8081444, 24'd8400969, 24'd8718048, 24'd8969931, 24'd9106771, 24'd9101488, 24'd8955127, 24'd8696653, 
24'd8377218, 24'd8060036, 24'd7807878, 24'd7670645, 24'd7675496, 24'd7821470, 24'd8079680, 24'd8399026, 24'd8716310, 24'd8968742, 24'd9106367, 24'd9101948, 24'd8956361, 24'd8698416, 24'd8379161, 24'd8061775, 24'd7809069, 24'd7671052, 24'd7675038, 24'd7820238, 24'd8077918, 24'd8397082, 24'd8714569, 24'd8967549, 24'd9105958, 24'd9102404, 24'd8957591, 24'd8700177, 24'd8381105, 24'd8063517, 
24'd7810264, 24'd7671464, 24'd7674585, 24'd7819011, 24'd8076158, 24'd8395139, 24'd8712827, 24'd8966352, 24'd9105544, 24'd9102854, 24'd8958817, 24'd8701936, 24'd8383048, 24'd8065260, 24'd7811462, 24'd7671880, 24'd7674137, 24'd7817787, 24'd8074400, 24'd8393195, 24'd8711082, 24'd8965152, 24'd9105124, 24'd9103300, 24'd8960039, 24'd8703693, 24'd8384992, 24'd8067006, 24'd7812665, 24'd7672302, 
24'd7673695, 24'd7816567, 24'd8072645, 24'd8391252, 24'd8709335, 24'd8963947, 24'd9104700, 24'd9103740, 24'd8961257, 24'd8705447, 24'd8386935, 24'd8068755, 24'd7813872, 24'd7672729, 24'd7673257, 24'd7815351, 24'd8070892, 24'd8389308, 24'd8707585, 24'd8962738, 24'd9104271, 24'd9104175, 24'd8962470, 24'd8707199, 24'd8388879, 24'd8070505, 24'd7815083, 24'd7673161, 24'd7672824, 24'd7814139, 
24'd8069141, 24'd8387364, 24'd8705834, 24'd8961525, 24'd9103837, 24'd9104606, 24'd8963680, 24'd8708949, 24'd8390822, 24'd8072258, 24'd7816298, 24'd7673597, 24'd7672396, 24'd7812931, 24'd8067392, 24'd8385421, 24'd8704080, 24'd8960308, 24'd9103397, 24'd9105031, 24'd8964886, 24'd8710696, 24'd8392766, 24'd8074013, 24'd7817517, 24'd7674039, 24'd7671973, 24'd7811728, 24'd8065646, 24'd8383477, 
24'd8702324, 24'd8959087, 24'd9102953, 24'd9105451, 24'd8966088, 24'd8712442, 24'd8394709, 24'd8075770, 24'd7818740, 24'd7674486, 24'd7671555, 24'd7810528, 24'd8063902, 24'd8381534, 24'd8700566, 24'd8957862, 24'd9102504, 24'd9105867, 24'd8967285, 24'd8714185, 24'd8396653, 24'd8077529, 24'd7819967, 24'd7674938, 24'd7671143, 24'd7809332, 24'd8062160, 24'd8379590, 24'd8698805, 24'd8956633, 
24'd9102049, 24'd9106277, 24'd8968479, 24'd8715925, 24'd8398596, 24'd8079291, 24'd7821198, 24'd7675395, 24'd7670735, 24'd7808141, 24'd8060420, 24'd8377647, 24'd8697043, 24'd8955400, 24'd9101590, 24'd9106682, 24'd8969669, 24'd8717664, 24'd8400540, 24'd8081054, 24'd7822433, 24'd7675856, 24'd7670332, 24'd7806953, 24'd8058683, 24'd8375704, 24'd8695278, 24'd8954163, 24'd9101126, 24'd9107082, 
24'd8970854, 24'd8719400, 24'd8402483, 24'd8082820, 24'd7823672, 24'd7676323, 24'd7669934, 24'd7805770, 24'd8056948, 24'd8373760, 24'd8693511, 24'd8952922, 24'd9100657, 24'd9107477, 24'd8972035, 24'd8721134, 24'd8404426, 24'd8084588, 24'd7824915, 24'd7676795, 24'd7669542, 24'd7804590, 24'd8055215, 24'd8371817, 24'd8691742, 24'd8951678, 24'd9100182, 24'd9107868, 24'd8973213, 24'd8722866, 
24'd8406369, 24'd8086358, 24'd7826161, 24'd7677272, 24'd7669154, 24'd7803415, 24'd8053485, 24'd8369874, 24'd8689971, 24'd8950429, 24'd9099703, 24'd9108253, 24'd8974386, 24'd8724595, 24'd8408312, 24'd8088130, 24'd7827412, 24'd7677754, 24'd7668772, 24'd7802244, 24'd8051757, 24'd8367931, 24'd8688198, 24'd8949176, 24'd9099219, 24'd9108633, 24'd8975555, 24'd8726322, 24'd8410255, 24'd8089905, 
24'd7828667, 24'd7678240, 24'd7668394, 24'd7801077, 24'd8050031, 24'd8365989, 24'd8686423, 24'd8947919, 24'd9098729, 24'd9109008, 24'd8976720, 24'd8728046, 24'd8412198, 24'd8091681, 24'd7829925, 24'd7678732, 24'd7668022, 24'd7799914, 24'd8048308, 24'd8364046, 24'd8684645, 24'd8946659, 24'd9098235, 24'd9109378, 24'd8977881, 24'd8729768, 24'd8414140, 24'd8093459, 24'd7831188, 24'd7679229, 
24'd7667654, 24'd7798755, 24'd8046587, 24'd8362104, 24'd8682866, 24'd8945394, 24'd9097736, 24'd9109742, 24'd8979038, 24'd8731488, 24'd8416082, 24'd8095240, 24'd7832454, 24'd7679730, 24'd7667292, 24'd7797601, 24'd8044868, 24'd8360161, 24'd8681084, 24'd8944126, 24'd9097232, 24'd9110102, 24'd8980190, 24'd8733205, 24'd8418025, 24'd8097023, 24'd7833725, 24'd7680237, 24'd7666935, 24'd7796450, 
24'd8043152, 24'd8358219, 24'd8679300, 24'd8942854, 24'd9096723, 24'd9110457, 24'd8981339, 24'd8734920, 24'd8419967, 24'd8098807, 24'd7834999, 24'd7680749, 24'd7666583, 24'd7795304, 24'd8041439, 24'd8356278, 24'd8677515, 24'd8941577, 24'd9096209, 24'd9110807, 24'd8982483, 24'd8736632, 24'd8421908, 24'd8100594, 24'd7836277, 24'd7681265, 24'd7666235, 24'd7794161, 24'd8039727, 24'd8354336, 
24'd8675727, 24'd8940297, 24'd9095689, 24'd9111151, 24'd8983623, 24'd8738342, 24'd8423850, 24'd8102383, 24'd7837559, 24'd7681787, 24'd7665893, 24'd7793023, 24'd8038019, 24'd8352395, 24'd8673937, 24'd8939014, 24'd9095165, 24'd9111491, 24'd8984759, 24'd8740050, 24'd8425791, 24'd8104173, 24'd7838845, 24'd7682313, 24'd7665556, 24'd7791890, 24'd8036312, 24'd8350454, 24'd8672146, 24'd8937726, 
24'd9094636, 24'd9111825, 24'd8985891, 24'd8741755, 24'd8427732, 24'd8105966, 24'd7840135, 24'd7682845, 24'd7665224, 24'd7790760, 24'd8034608, 24'd8348513, 24'd8670352, 24'd8936434, 24'd9094103, 24'd9112155, 24'd8987018, 24'd8743458, 24'd8429673, 24'd8107761, 24'd7841428, 24'd7683381, 24'd7664897, 24'd7789634, 24'd8032907, 24'd8346572, 24'd8668556, 24'd8935139, 24'd9093564, 24'd9112479, 
24'd8988142, 24'd8745158, 24'd8431613, 24'd8109557, 24'd7842726, 24'd7683923, 24'd7664576, 24'd7788513, 24'd8031208, 24'd8344632, 24'd8666758, 24'd8933839, 24'd9093020, 24'd9112798, 24'd8989261, 24'd8746855, 24'd8433553, 24'd8111356, 24'd7844027, 24'd7684469, 24'd7664259, 24'd7787396, 24'd8029512, 24'd8342692, 24'd8664959, 24'd8932536, 24'd9092471, 24'd9113113, 24'd8990376, 24'd8748550, 
24'd8435493, 24'd8113157, 24'd7845332, 24'd7685020, 24'd7663947, 24'd7786283, 24'd8027818, 24'd8340752, 24'd8663157, 24'd8931229, 24'd9091917, 24'd9113422, 24'd8991487, 24'd8750243, 24'd8437432, 24'd8114959, 24'd7846641, 24'd7685576, 24'd7663641, 24'd7785175, 24'd8026127, 24'd8338813, 24'd8661354, 24'd8929919, 24'd9091359, 24'd9113726, 24'd8992593, 24'd8751933, 24'd8439371, 24'd8116764, 
24'd7847953, 24'd7686137, 24'd7663339, 24'd7784070, 24'd8024438, 24'd8336874, 24'd8659549, 24'd8928604, 24'd9090795, 24'd9114025, 24'd8993695, 24'd8753620, 24'd8441310, 24'd8118570, 24'd7849270, 24'd7686703, 24'd7663043, 24'd7782970, 24'd8022752, 24'd8334936, 24'd8657741, 24'd8927286, 24'd9090227, 24'd9114319, 24'd8994794, 24'd8755305, 24'd8443248, 24'd8120378, 24'd7850590, 24'd7687274, 
24'd7662751, 24'd7781874, 24'd8021068, 24'd8332998, 24'd8655932, 24'd8925964, 24'd9089653, 24'd9114607, 24'd8995887, 24'd8756988, 24'd8445186, 24'd8122188, 24'd7851914, 24'd7687850, 24'd7662465, 24'd7780782, 24'd8019387, 24'd8331060, 24'd8654121, 24'd8924638, 24'd9089075, 24'd9114891, 24'd8996977, 24'd8758668, 24'd8447124, 24'd8124000, 24'd7853242, 24'd7688431, 24'd7662184, 24'd7779695, 
24'd8017709, 24'd8329122, 24'd8652308, 24'd8923308, 24'd9088492, 24'd9115170, 24'd8998062, 24'd8760345, 24'd8449061, 24'd8125814, 24'd7854573, 24'd7689017, 24'd7661908, 24'd7778612, 24'd8016033, 24'd8327185, 24'd8650493, 24'd8921975, 24'd9087904, 24'd9115443, 24'd8999143, 24'd8762019, 24'd8450998, 24'd8127630, 24'd7855908, 24'd7689607, 24'd7661637, 24'd7777533, 24'd8014359, 24'd8325249, 
24'd8648677, 24'd8920638, 24'd9087311, 24'd9115712, 24'd9000220, 24'd8763691, 24'd8452934, 24'd8129447, 24'd7857247, 24'd7690203, 24'd7661371, 24'd7776458, 24'd8012689, 24'd8323313, 24'd8646858, 24'd8919297, 24'd9086713, 24'd9115975, 24'd9001292, 24'd8765361, 24'd8454870, 24'd8131266, 24'd7858590, 24'd7690803, 24'd7661110, 24'd7775388, 24'd8011021, 24'd8321377, 24'd8645038, 24'd8917952, 
24'd9086110, 24'd9116233, 24'd9002360, 24'd8767027, 24'd8456806, 24'd8133088, 24'd7859936, 24'd7691408, 24'd7660855, 24'd7774322, 24'd8009355, 24'd8319442, 24'd8643216, 24'd8916604, 24'd9085502, 24'd9116486, 24'd9003424, 24'd8768691, 24'd8458740, 24'd8134910, 24'd7861287, 24'd7692019, 24'd7660604, 24'd7773260, 24'd8007693, 24'd8317507, 24'd8641392, 24'd8915252, 24'd9084890, 24'd9116734, 
24'd9004484, 24'd8770353, 24'd8460675, 24'd8136735, 24'd7862640, 24'd7692634, 24'd7660359, 24'd7772203, 24'd8006033, 24'd8315573, 24'd8639567, 24'd8913896, 24'd9084272, 24'd9116977, 24'd9005539, 24'd8772011, 24'd8462609, 24'd8138562, 24'd7863998, 24'd7693254, 24'd7660118, 24'd7771150, 24'd8004375, 24'd8313639, 24'd8637740, 24'd8912537, 24'd9083650, 24'd9117215, 24'd9006590, 24'd8773667, 
24'd8464542, 24'd8140390, 24'd7865359, 24'd7693878, 24'd7659883, 24'd7770101, 24'd8002721, 24'd8311706, 24'd8635911, 24'd8911174, 24'd9083022, 24'd9117448, 24'd9007636, 24'd8775321, 24'd8466475, 24'd8142220, 24'd7866724, 24'd7694508, 24'd7659653, 24'd7769057, 24'd8001069, 24'd8309774, 24'd8634080, 24'd8909807, 24'd9082390, 24'd9117675, 24'd9008679, 24'd8776971, 24'd8468407, 24'd8144051, 
24'd7868092, 24'd7695143, 24'd7659428, 24'd7768017, 24'd7999419, 24'd8307842, 24'd8632247, 24'd8908437, 24'd9081753, 24'd9117898, 24'd9009717, 24'd8778619, 24'd8470339, 24'd8145885, 24'd7869465, 24'd7695782, 24'd7659208, 24'd7766981, 24'd7997773, 24'd8305910, 24'd8630413, 24'd8907063, 24'd9081112, 24'd9118115, 24'd9010750, 24'd8780264, 24'd8472270, 24'd8147720, 24'd7870840, 24'd7696426, 
24'd7658993, 24'd7765950, 24'd7996129, 24'd8303979, 24'd8628577, 24'd8905685, 24'd9080465, 24'd9118327, 24'd9011779, 24'd8781907, 24'd8474201, 24'd8149557, 24'd7872220, 24'd7697075, 24'd7658784, 24'd7764923, 24'd7994488, 24'd8302049, 24'd8626739, 24'd8904304, 24'd9079813, 24'd9118534, 24'd9012804, 24'd8783546, 24'd8476131, 24'd8151395, 24'd7873603, 24'd7697729, 24'd7658579, 24'd7763900, 
24'd7992850, 24'd8300119, 24'd8624900, 24'd8902919, 24'd9079157, 24'd9118736, 24'd9013824, 24'd8785183, 24'd8478060, 24'd8153235, 24'd7874990, 24'd7698388, 24'd7658380, 24'd7762882, 24'd7991214, 24'd8298190, 24'd8623059, 24'd8901531, 24'd9078496, 24'd9118933, 24'd9014840, 24'd8786817, 24'd8479989, 24'd8155077, 24'd7876380, 24'd7699052, 24'd7658185, 24'd7761868, 24'd7989582, 24'd8296262, 
24'd8621217, 24'd8900139, 24'd9077830, 24'd9119125, 24'd9015852, 24'd8788449, 24'd8481917, 24'd8156920, 24'd7877774, 24'd7699720, 24'd7657996, 24'd7760859, 24'd7987952, 24'd8294334, 24'd8619372, 24'd8898743, 24'd9077159, 24'd9119311, 24'd9016859, 24'd8790077, 24'd8483845, 24'd8158765, 24'd7879171, 24'd7700393, 24'd7657812, 24'd7759854, 24'd7986325, 24'd8292407, 24'd8617527, 24'd8897344, 
24'd9076483, 24'd9119493, 24'd9017862, 24'd8791703, 24'd8485772, 24'd8160612, 24'd7880572, 24'd7701072, 24'd7657633, 24'd7758853, 24'd7984700, 24'd8290480, 24'd8615679, 24'd8895941, 24'd9075802, 24'd9119669, 24'd9018860, 24'd8793326, 24'd8487698, 24'd8162460, 24'd7881977, 24'd7701755, 24'd7657459, 24'd7757857, 24'd7983079, 24'd8288554, 24'd8613830, 24'd8894535, 24'd9075117, 24'd9119841, 
24'd9019854, 24'd8794946, 24'd8489623, 24'd8164310, 24'd7883385, 24'd7702442, 24'd7657291, 24'd7756865, 24'd7981460, 24'd8286629, 24'd8611979, 24'd8893125, 24'd9074427, 24'd9120007, 24'd9020844, 24'd8796563, 24'd8491548, 24'd8166161, 24'd7884797, 24'd7703135, 24'd7657127, 24'd7755878, 24'd7979845, 24'd8284705, 24'd8610127, 24'd8891711, 24'd9073732, 24'd9120168, 24'd9021829, 24'd8798177, 
24'd8493472, 24'd8168014, 24'd7886212, 24'd7703832, 24'd7656969, 24'd7754895, 24'd7978232, 24'd8282781, 24'd8608274, 24'd8890294, 24'd9073032, 24'd9120324, 24'd9022810, 24'd8799789, 24'd8495395, 24'd8169869, 24'd7887630, 24'd7704535, 24'd7656815, 24'd7753917, 24'd7976622, 24'd8280858, 24'd8606418, 24'd8888874, 24'd9072328, 24'd9120474, 24'd9023786, 24'd8801397, 24'd8497318, 24'd8171725, 
24'd7889053, 24'd7705242, 24'd7656667, 24'd7752942, 24'd7975015, 24'd8278936, 24'd8604562, 24'd8887450, 24'd9071618, 24'd9120620, 24'd9024758, 24'd8803003, 24'd8499240, 24'd8173582, 24'd7890478, 24'd7705953, 24'd7656524, 24'd7751973, 24'd7973411, 24'd8277015, 24'd8602703, 24'd8886022, 24'd9070904, 24'd9120760, 24'd9025725, 24'd8804605, 24'd8501161, 24'd8175442, 24'd7891908, 24'd7706670, 
24'd7656386, 24'd7751008, 24'd7971809, 24'd8275094, 24'd8600843, 24'd8884591, 24'd9070185, 24'd9120896, 24'd9026688, 24'd8806205, 24'd8503081, 24'd8177302, 24'd7893340, 24'd7707391, 24'd7656253, 24'd7750047, 24'd7970211, 24'd8273174, 24'd8598982, 24'd8883157, 24'd9069461, 24'd9121026, 24'd9027646, 24'd8807802, 24'd8505000, 24'd8179164, 24'd7894777, 24'd7708117, 24'd7656126, 24'd7749091, 
24'd7968615, 24'd8271256, 24'd8597119, 24'd8881719, 24'd9068733, 24'd9121151, 24'd9028600, 24'd8809396, 24'd8506919, 24'd8181028, 24'd7896216, 24'd7708848, 24'd7656003, 24'd7748139, 24'd7967023, 24'd8269337, 24'd8595255, 24'd8880278, 24'd9068000, 24'd9121271, 24'd9029550, 24'd8810987, 24'd8508836, 24'd8182893, 24'd7897659, 24'd7709584, 24'd7655886, 24'd7747192, 24'd7965433, 24'd8267420, 
24'd8593389, 24'd8878833, 24'd9067262, 24'd9121386, 24'd9030495, 24'd8812575, 24'd8510753, 24'd8184759, 24'd7899106, 24'd7710324, 24'd7655774, 24'd7746250, 24'd7963847, 24'd8265504, 24'd8591522, 24'd8877385, 24'd9066519, 24'd9121496, 24'd9031435, 24'd8814160, 24'd8512669, 24'd8186627, 24'd7900556, 24'd7711069, 24'd7655667, 24'd7745311, 24'd7962263, 24'd8263588, 24'd8589654, 24'd8875933, 
24'd9065771, 24'd9121600, 24'd9032371, 24'd8815742, 24'd8514585, 24'd8188496, 24'd7902009, 24'd7711819, 24'd7655565, 24'd7744378, 24'd7960683, 24'd8261673, 24'd8587784, 24'd8874478, 24'd9065019, 24'd9121699, 24'd9033302, 24'd8817321, 24'd8516499, 24'd8190367, 24'd7903466, 24'd7712574, 24'd7655468, 24'd7743449, 24'd7959105, 24'd8259759, 24'd8585912, 24'd8873019, 24'd9064262, 24'd9121794, 
24'd9034229, 24'd8818898, 24'd8518412, 24'd8192239, 24'd7904926, 24'd7713333, 24'd7655376, 24'd7742524, 24'd7957530, 24'd8257846, 24'd8584040, 24'd8871557, 24'd9063500, 24'd9121883, 24'd9035152, 24'd8820471, 24'd8520325, 24'd8194112, 24'd7906390, 24'd7714098, 24'd7655290, 24'd7741604, 24'd7955959, 24'd8255934, 24'd8582166, 24'd8870092, 24'd9062734, 24'd9121967, 24'd9036070, 24'd8822041, 
24'd8522236, 24'd8195987, 24'd7907857, 24'd7714866, 24'd7655208, 24'd7740688, 24'd7954390, 24'd8254023, 24'd8580290, 24'd8868623, 24'd9061962, 24'd9122046, 24'd9036983, 24'd8823608, 24'd8524147, 24'd8197863, 24'd7909327, 24'd7715640, 24'd7655132, 24'd7739777, 24'd7952825, 24'd8252113, 24'd8578413, 24'd8867151, 24'd9061186, 24'd9122119, 24'd9037892, 24'd8825172, 24'd8526057, 24'd8199741, 
24'd7910801, 24'd7716418, 24'd7655061, 24'd7738871, 24'd7951262, 24'd8250204, 24'd8576535, 24'd8865676, 24'd9060406, 24'd9122188, 24'd9038796, 24'd8826733, 24'd8527965, 24'd8201619, 24'd7912278, 24'd7717201, 24'd7654995, 24'd7737969, 24'd7949703, 24'd8248296, 24'd8574656, 24'd8864197, 24'd9059620, 24'd9122251, 24'd9039695, 24'd8828290, 24'd8529873, 24'd8203499, 24'd7913758, 24'd7717989, 
24'd7654934, 24'd7737072, 24'd7948147, 24'd8246388, 24'd8572775, 24'd8862715, 24'd9058830, 24'd9122309, 24'd9040590, 24'd8829845, 24'd8531780, 24'd8205381, 24'd7915242, 24'd7718782, 24'd7654878, 24'd7736179, 24'd7946594, 24'd8244482, 24'd8570893, 24'd8861230, 24'd9058035, 24'd9122363, 24'd9041481, 24'd8831397, 24'd8533686, 24'd8207264, 24'd7916729, 24'd7719579, 24'd7654828, 24'd7735291, 
24'd7945044, 24'd8242577, 24'd8569010, 24'd8859741, 24'd9057236, 24'd9122411, 24'd9042367, 24'd8832945, 24'd8535590, 24'd8209148, 24'd7918220, 24'd7720381, 24'd7654782, 24'd7734407, 24'd7943497, 24'd8240673, 24'd8567125, 24'd8858249, 24'd9056432, 24'd9122453, 24'd9043248, 24'd8834491, 24'd8537494, 24'd8211033, 24'd7919713, 24'd7721187, 24'd7654742, 24'd7733528, 24'd7941953, 24'd8238770, 
24'd8565239, 24'd8856754, 24'd9055623, 24'd9122491, 24'd9044125, 24'd8836033, 24'd8539397, 24'd8212919, 24'd7921210, 24'd7721998, 24'd7654707, 24'd7732653, 24'd7940412, 24'd8236867, 24'd8563352, 24'd8855255, 24'd9054809, 24'd9122524, 24'd9044997, 24'd8837572, 24'd8541298, 24'd8214807, 24'd7922710, 24'd7722814, 24'd7654677, 24'd7731784, 24'd7938874, 24'd8234966, 24'd8561464, 24'd8853753, 
24'd9053991, 24'd9122551, 24'd9045865, 24'd8839108, 24'd8543199, 24'd8216696, 24'd7924214, 24'd7723635, 24'd7654652, 24'd7730918, 24'd7937340, 24'd8233066, 24'd8559574, 24'd8852248, 24'd9053168, 24'd9122573, 24'd9046728, 24'd8840641, 24'd8545098, 24'd8218586, 24'd7925721, 24'd7724460, 24'd7654633, 24'd7730058, 24'd7935809, 24'd8231168, 24'd8557684, 24'd8850740, 24'd9052341, 24'd9122590, 
24'd9047586, 24'd8842171, 24'd8546996, 24'd8220477, 24'd7927231, 24'd7725290, 24'd7654618, 24'd7729202, 24'd7934281, 24'd8229270, 24'd8555792, 24'd8849228, 24'd9051509, 24'd9122602, 24'd9048440, 24'd8843697, 24'd8548894, 24'd8222370, 24'd7928744, 24'd7726124, 24'd7654609, 24'd7728350, 24'd7932756, 24'd8227373, 24'd8553899, 24'd8847713, 24'd9050672, 24'd9122609, 24'd9049289, 24'd8845221, 
24'd8550790, 24'd8224263, 24'd7930260, 24'd7726963, 24'd7654605, 24'd7727504, 24'd7931234, 24'd8225478, 24'd8552004, 24'd8846195, 24'd9049830, 24'd9122611, 24'd9050133, 24'd8846741, 24'd8552685, 24'd8226158, 24'd7931780, 24'd7727807, 24'd7654605, 24'd7726661, 24'd7929715, 24'd8223583, 24'd8550109, 24'd8844674, 24'd9048984, 24'd9122607, 24'd9050973, 24'd8848258, 24'd8554579, 24'd8228054, 
24'd7933303, 24'd7728656, 24'd7654612, 24'd7725824, 24'd7928200, 24'd8221690, 24'd8548212, 24'd8843149, 24'd9048133, 24'd9122598, 24'd9051808, 24'd8849771, 24'd8556471, 24'd8229951, 24'd7934829, 24'd7729509, 24'd7654623, 24'd7724991, 24'd7926688, 24'd8219798, 24'd8546315, 24'd8841622, 24'd9047278, 24'd9122585, 24'd9052639, 24'd8851282, 24'd8558363, 24'd8231849, 24'd7936358, 24'd7730366, 
24'd7654639, 24'd7724163, 24'd7925179, 24'd8217907, 24'd8544416, 24'd8840091, 24'd9046418, 24'd9122566, 24'd9053464, 24'd8852789, 24'd8560253, 24'd8233749, 24'd7937891, 24'd7731229, 24'd7654661, 24'd7723339, 24'd7923674, 24'd8216017, 24'd8542516, 24'd8838557, 24'd9045554, 24'd9122542, 24'd9054286, 24'd8854293, 24'd8562142, 24'd8235649, 24'd7939426, 24'd7732095, 24'd7654687, 24'd7722521, 
24'd7922171, 24'd8214129, 24'd8540615, 24'd8837020, 24'd9044684, 24'd9122512, 24'd9055102, 24'd8855794, 24'd8564030, 24'd8237550, 24'd7940965, 24'd7732967, 24'd7654719, 24'd7721706, 24'd7920672, 24'd8212242, 24'd8538713, 24'd8835480, 24'd9043811, 24'd9122478, 24'd9055914, 24'd8857291, 24'd8565917, 24'd8239453, 24'd7942507, 24'd7733843, 24'd7654756, 24'd7720897, 24'd7919176, 24'd8210356, 
24'd8536810, 24'd8833936, 24'd9042932, 24'd9122439, 24'd9056721, 24'd8858785, 24'd8567802, 24'd8241357, 24'd7944052, 24'd7734724, 24'd7654798, 24'd7720092, 24'd7917684, 24'd8208471, 24'd8534906, 24'd8832390, 24'd9042049, 24'd9122394, 24'd9057524, 24'd8860276, 24'd8569686, 24'd8243261, 24'd7945600, 24'd7735609, 24'd7654845, 24'd7719292, 24'd7916195, 24'd8206587, 24'd8533001, 24'd8830840, 
24'd9041162, 24'd9122344, 24'd9058321, 24'd8861764, 24'd8571569, 24'd8245167, 24'd7947151, 24'd7736499, 24'd7654898, 24'd7718496, 24'd7914709, 24'd8204705, 24'd8531095, 24'd8829287, 24'd9040269, 24'd9122289, 24'd9059114, 24'd8863248, 24'd8573451, 24'd8247073, 24'd7948705, 24'd7737393, 24'd7654955, 24'd7717706, 24'd7913226, 24'd8202824, 24'd8529188, 24'd8827731, 24'd9039373, 24'd9122229, 
24'd9059903, 24'd8864729, 24'd8575331, 24'd8248981, 24'd7950263, 24'd7738292, 24'd7655018, 24'd7716920, 24'd7911747, 24'd8200944, 24'd8527280, 24'd8826172, 24'd9038472, 24'd9122164, 24'd9060687, 24'd8866206, 24'd8577210, 24'd8250890, 24'd7951823, 24'd7739196, 24'd7655086, 24'd7716138, 24'd7910271, 24'd8199066, 24'd8525371, 24'd8824610, 24'd9037566, 24'd9122093, 24'd9061466, 24'd8867680, 
24'd8579088, 24'd8252799, 24'd7953387, 24'd7740104, 24'd7655159, 24'd7715362, 24'd7908799, 24'd8197189, 24'd8523461, 24'd8823045, 24'd9036655, 24'd9122018, 24'd9062240, 24'd8869151, 24'd8580964, 24'd8254710, 24'd7954953, 24'd7741017, 24'd7655237, 24'd7714590, 24'd7907330, 24'd8195313, 24'd8521550, 24'd8821477, 24'd9035740, 24'd9121937, 24'd9063009, 24'd8870619, 24'd8582839, 24'd8256621, 
24'd7956523, 24'd7741934, 24'd7655320, 24'd7713823, 24'd7905864, 24'd8193439, 24'd8519638, 24'd8819906, 24'd9034821, 24'd9121851, 24'd9063774, 24'd8872083, 24'd8584712, 24'd8258533, 24'd7958096, 24'd7742855, 24'd7655408, 24'd7713060, 24'd7904401, 24'd8191566, 24'd8517725, 24'd8818332, 24'd9033897, 24'd9121760, 24'd9064534, 24'd8873543, 24'd8586585, 24'd8260447, 24'd7959671, 24'd7743782, 
24'd7655502, 24'd7712302, 24'd7902942, 24'd8189695, 24'd8515811, 24'd8816755, 24'd9032968, 24'd9121664, 24'd9065290, 24'd8875001, 24'd8588456, 24'd8262361, 24'd7961250, 24'd7744712, 24'd7655601, 24'd7711550, 24'd7901487, 24'd8187825, 24'd8513897, 24'd8815175, 24'd9032035, 24'd9121563, 24'd9066040, 24'd8876455, 24'd8590325, 24'd8264276, 24'd7962832, 24'd7745648, 24'd7655704, 24'd7710801, 
24'd7900035, 24'd8185956, 24'd8511981, 24'd8813591, 24'd9031098, 24'd9121457, 24'd9066786, 24'd8877905, 24'd8592193, 24'd8266192, 24'd7964416, 24'd7746588, 24'd7655813, 24'd7710058, 24'd7898586, 24'd8184089, 24'd8510065, 24'd8812005, 24'd9030156, 24'd9121345, 24'd9067527, 24'd8879352, 24'd8594060, 24'd8268109, 24'd7966004, 24'd7747532, 24'd7655927, 24'd7709319, 24'd7897141, 24'd8182223, 
24'd8508148, 24'd8810416, 24'd9029209, 24'd9121229, 24'd9068263, 24'd8880796, 24'd8595925, 24'd8270026, 24'd7967595, 24'd7748481, 24'd7656047, 24'd7708585, 24'd7895699, 24'd8180358, 24'd8506230, 24'd8808824, 24'd9028258, 24'd9121107, 24'd9068995, 24'd8882236, 24'd8597788, 24'd8271945, 24'd7969188, 24'd7749434, 24'd7656171, 24'd7707856, 24'd7894260, 24'd8178495, 24'd8504311, 24'd8807229, 
24'd9027303, 24'd9120980, 24'd9069722, 24'd8883673, 24'd8599651, 24'd8273864, 24'd7970785, 24'd7750392, 24'd7656301, 24'd7707132, 24'd7892825, 24'd8176634, 24'd8502391, 24'd8805631, 24'd9026343, 24'd9120848, 24'd9070444, 24'd8885106, 24'd8601512, 24'd8275784, 24'd7972384, 24'd7751354, 24'd7656435, 24'd7706412, 24'd7891394, 24'd8174774, 24'd8500471, 24'd8804030, 24'd9025378, 24'd9120711, 
24'd9071161, 24'd8886535, 24'd8603371, 24'd8277705, 24'd7973986, 24'd7752321, 24'd7656575, 24'd7705697, 24'd7889966, 24'd8172915, 24'd8498549, 24'd8802426, 24'd9024409, 24'd9120568, 24'd9071874, 24'd8887962, 24'd8605229, 24'd8279627, 24'd7975592, 24'd7753292, 24'd7656720, 24'd7704987, 24'd7888542, 24'd8171058, 24'd8496627, 24'd8800820, 24'd9023436, 24'd9120421, 24'd9072581, 24'd8889384, 
24'd8607085, 24'd8281549, 24'd7977200, 24'd7754267, 24'd7656870, 24'd7704282, 24'd7887121, 24'd8169203, 24'd8494705, 24'd8799210, 24'd9022458, 24'd9120268, 24'd9073284, 24'd8890804, 24'd8608940, 24'd8283472, 24'd7978811, 24'd7755247, 24'd7657025, 24'd7703581, 24'd7885703, 24'd8167349, 24'd8492781, 24'd8797598, 24'd9021476, 24'd9120111, 24'd9073982, 24'd8892219, 24'd8610793, 24'd8285396, 
24'd7980425, 24'd7756232, 24'd7657185, 24'd7702886, 24'd7884289, 24'd8165496, 24'd8490857, 24'd8795982, 24'd9020489, 24'd9119948, 24'd9074675, 24'd8893631, 24'd8612644, 24'd8287321, 24'd7982041, 24'd7757221, 24'd7657351, 24'd7702195, 24'd7882879, 24'd8163645, 24'd8488932, 24'd8794364, 24'd9019498, 24'd9119780, 24'd9075364, 24'd8895040, 24'd8614494, 24'd8289246, 24'd7983661, 24'd7758214, 
24'd7657521, 24'd7701509, 24'd7881472, 24'd8161796, 24'd8487006, 24'd8792743, 24'd9018502, 24'd9119607, 24'd9076047, 24'd8896445, 24'd8616343, 24'd8291172, 24'd7985283, 24'd7759212, 24'd7657697, 24'd7700828, 24'd7880069, 24'd8159949, 24'd8485080, 24'd8791119, 24'd9017502, 24'd9119428, 24'd9076726, 24'd8897847, 24'd8618190, 24'd8293099, 24'd7986909, 24'd7760214, 24'd7657878, 24'd7700151, 
24'd7878669, 24'd8158103, 24'd8483153, 24'd8789493, 24'd9016498, 24'd9119245, 24'd9077400, 24'd8899245, 24'd8620035, 24'd8295026, 24'd7988537, 24'd7761221, 24'd7658064, 24'd7699480, 24'd7877273, 24'd8156258, 24'd8481225, 24'd8787863, 24'd9015489, 24'd9119057, 24'd9078069, 24'd8900639, 24'd8621879, 24'd8296954, 24'd7990168, 24'd7762232, 24'd7658255, 24'd7698813, 24'd7875880, 24'd8154415, 
24'd8479297, 24'd8786231, 24'd9014476, 24'd9118863, 24'd9078734, 24'd8902030, 24'd8623721, 24'd8298883, 24'd7991801, 24'd7763247, 24'd7658451, 24'd7698151, 24'd7874491, 24'd8152574, 24'd8477368, 24'd8784596, 24'd9013458, 24'd9118664, 24'd9079393, 24'd8903417, 24'd8625561, 24'd8300812, 24'd7993438, 24'd7764267, 24'd7658652, 24'd7697494, 24'd7873106, 24'd8150735, 24'd8475438, 24'd8782958, 
24'd9012436, 24'd9118460, 24'd9080048, 24'd8904801, 24'd8627400, 24'd8302742, 24'd7995077, 24'd7765291, 24'd7658858, 24'd7696842, 24'd7871724, 24'd8148897, 24'd8473508, 24'd8781317, 24'd9011410, 24'd9118251, 24'd9080698, 24'd8906180, 24'd8629237, 24'd8304673, 24'd7996719, 24'd7766320, 24'd7659070, 24'd7696194, 24'd7870346, 24'd8147061, 24'd8471577, 24'd8779674, 24'd9010379, 24'd9118037, 
24'd9081343, 24'd8907557, 24'd8631072, 24'd8306604, 24'd7998364, 24'd7767353, 24'd7659287, 24'd7695552, 24'd7868971, 24'd8145226, 24'd8469646, 24'd8778028, 24'd9009344, 24'd9117818, 24'd9081983, 24'd8908929, 24'd8632906, 24'd8308535, 24'd8000011, 24'd7768390, 24'd7659508, 24'd7694914, 24'd7867601, 24'd8143393, 24'd8467714, 24'd8776379, 24'd9008305, 24'd9117594, 24'd9082618, 24'd8910299, 
24'd8634737, 24'd8310468, 24'd8001662, 24'd7769431, 24'd7659735, 24'd7694281, 24'd7866233, 24'd8141562, 24'd8465781, 24'd8774727, 24'd9007261, 24'd9117365, 24'd9083248, 24'd8911664, 24'd8636568, 24'd8312400, 24'd8003315, 24'd7770477, 24'd7659967, 24'd7693653, 24'd7864870, 24'd8139733, 24'd8463848, 24'd8773073, 24'd9006213, 24'd9117130, 24'd9083874, 24'd8913026, 24'd8638396, 24'd8314334, 
24'd8004970, 24'd7771528, 24'd7660204, 24'd7693030, 24'd7863510, 24'd8137905, 24'd8461914, 24'd8771416, 24'd9005161, 24'd9116890, 24'd9084494, 24'd8914384, 24'd8640223, 24'd8316268, 24'd8006629, 24'd7772582, 24'd7660446, 24'd7692412, 24'd7862154, 24'd8136080, 24'd8459980, 24'd8769756, 24'd9004104, 24'd9116646, 24'd9085110, 24'd8915738, 24'd8642048, 24'd8318202, 24'd8008289, 24'd7773641, 
24'd7660694, 24'd7691799, 24'd7860801, 24'd8134256, 24'd8458046, 24'd8768094, 24'd9003043, 24'd9116396, 24'd9085721, 24'd8917089, 24'd8643871, 24'd8320137, 24'd8009953, 24'd7774704, 24'd7660946, 24'd7691190, 24'd7859452, 24'd8132433, 24'd8456110, 24'd8766429, 24'd9001977, 24'd9116141, 24'd9086327, 24'd8918436, 24'd8645692, 24'd8322072, 24'd8011619, 24'd7775772, 24'd7661203, 24'd7690587, 
24'd7858107, 24'd8130613, 24'd8454175, 24'd8764761, 24'd9000908, 24'd9115881, 24'd9086928, 24'd8919779, 24'd8647512, 24'd8324008, 24'd8013288, 24'd7776844, 24'd7661466, 24'd7689988, 24'd7856766, 24'd8128794, 24'd8452239, 24'd8763091, 24'd8999834, 24'd9115616, 24'd9087524, 24'd8921118, 24'd8649330, 24'd8325944, 24'd8014960, 24'd7777920, 24'd7661734, 24'd7689395, 24'd7855428, 24'd8126977, 
24'd8450302, 24'd8761418, 24'd8998755, 24'd9115345, 24'd9088115, 24'd8922454, 24'd8651145, 24'd8327881, 24'd8016634, 24'd7779000, 24'd7662007, 24'd7688806, 24'd7854094, 24'd8125162, 24'd8448365, 24'd8759743, 24'd8997673, 24'd9115070, 24'd9088702, 24'd8923786, 24'd8652959, 24'd8329818, 24'd8018311, 24'd7780085, 24'd7662284, 24'd7688222, 24'd7852764, 24'd8123349, 24'd8446428, 24'd8758065, 
24'd8996586, 24'd9114790, 24'd9089283, 24'd8925114, 24'd8654772, 24'd8331756, 24'd8019990, 24'd7781174, 24'd7662567, 24'd7687643, 24'd7851438, 24'd8121538, 24'd8444490, 24'd8756384, 24'd8995495, 24'd9114504, 24'd9089860, 24'd8926439, 24'd8656582, 24'd8333694, 24'd8021672, 24'd7782267, 24'd7662855, 24'd7687069, 24'd7850115, 24'd8119728, 24'd8442552, 24'd8754701, 24'd8994400, 24'd9114214, 
24'd9090431, 24'd8927760, 24'd8658391, 24'd8335632, 24'd8023357, 24'd7783365, 24'd7663149, 24'd7686500, 24'd7848796, 24'd8117921, 24'd8440614, 24'd8753015, 24'd8993300, 24'd9113918, 24'd9090998, 24'd8929077, 24'd8660197, 24'd8337571, 24'd8025044, 24'd7784466, 24'd7663447, 24'd7685935, 24'd7847481, 24'd8116115, 24'd8438675, 24'd8751326, 24'd8992196, 24'd9113617, 24'd9091560, 24'd8930390, 
24'd8662002, 24'd8339510, 24'd8026734, 24'd7785572, 24'd7663750, 24'd7685376, 24'd7846170, 24'd8114312, 24'd8436736, 24'd8749635, 24'd8991088, 24'd9113311, 24'd9092117, 24'd8931699, 24'd8663805, 24'd8341449, 24'd8028426, 24'd7786682, 24'd7664059, 24'd7684822, 24'd7844863, 24'd8112510, 24'd8434796, 24'd8747942, 24'd8989976, 24'd9113000, 24'd9092669, 24'd8933005, 24'd8665605, 24'd8343389, 
24'd8030121, 24'd7787797, 24'd7664372, 24'd7684272, 24'd7843559, 24'd8110710, 24'd8432856, 24'd8746246, 24'd8988859, 24'd9112684, 24'd9093216, 24'd8934306, 24'd8667404, 24'd8345329, 24'd8031818, 24'd7788915, 24'd7664691, 24'd7683728, 24'd7842259, 24'd8108912, 24'd8430916, 24'd8744547, 24'd8987739, 24'd9112363, 24'd9093758, 24'd8935604, 24'd8669201, 24'd8347269, 24'd8033518, 24'd7790038, 
24'd7665014, 24'd7683188, 24'd7840963, 24'd8107116, 24'd8428976, 24'd8742846, 24'd8986614, 24'd9112037, 24'd9094295, 24'd8936898, 24'd8670996, 24'd8349210, 24'd8035220, 24'd7791165, 24'd7665343, 24'd7682653, 24'd7839671, 24'd8105322, 24'd8427035, 24'd8741143, 24'd8985485, 24'd9111706, 24'd9094827, 24'd8938189, 24'd8672789, 24'd8351151, 24'd8036925, 24'd7792296, 24'd7665677, 24'd7682124, 
24'd7838383, 24'd8103530, 24'd8425094, 24'd8739437, 24'd8984352, 24'd9111370, 24'd9095354, 24'd8939475, 24'd8674580, 24'd8353092, 24'd8038632, 24'd7793432, 24'd7666016, 24'd7681599, 24'd7837098, 24'd8101740, 24'd8423152, 24'd8737728, 24'd8983214, 24'd9111028, 24'd9095876, 24'd8940758, 24'd8676369, 24'd8355033, 24'd8040342, 24'd7794571, 24'd7666359, 24'd7681079, 24'd7835818, 24'd8099952, 
24'd8421211, 24'd8736018, 24'd8982072, 24'd9110682, 24'd9096394, 24'd8942036, 24'd8678156, 24'd8356975, 24'd8042054, 24'd7795715, 24'd7666708, 24'd7680564, 24'd7834541, 24'd8098166, 24'd8419269, 24'd8734304, 24'd8980927, 24'd9110330, 24'd9096906, 24'd8943311, 24'd8679941, 24'd8358917, 24'd8043768, 24'd7796863, 24'd7667062, 24'd7680055, 24'd7833268, 24'd8096382, 24'd8417327, 24'd8732589, 
24'd8979777, 24'd9109974, 24'd9097413, 24'd8944582, 24'd8681724, 24'd8360859, 24'd8045485, 24'd7798015, 24'd7667422, 24'd7679550, 24'd7831999, 24'd8094600, 24'd8415385, 24'd8730870, 24'd8978623, 24'd9109612, 24'd9097916, 24'd8945849, 24'd8683505, 24'd8362801, 24'd8047205, 24'd7799171, 24'd7667786, 24'd7679050, 24'd7830734, 24'd8092820, 24'd8413443, 24'd8729150, 24'd8977464, 24'd9109245, 
24'd9098413, 24'd8947112, 24'd8685284, 24'd8364744, 24'd8048926, 24'd7800331, 24'd7668155, 24'd7678555, 24'd7829473, 24'd8091043, 24'd8411500, 24'd8727427, 24'd8976302, 24'd9108874, 24'd9098906, 24'd8948371, 24'd8687060, 24'd8366686, 24'd8050650, 24'd7801496, 24'd7668529, 24'd7678065, 24'd7828216, 24'd8089267, 24'd8409557, 24'd8725702, 24'd8975136, 24'd9108497, 24'd9099393, 24'd8949626, 
24'd8688835, 24'd8368629, 24'd8052377, 24'd7802664, 24'd7668909, 24'd7677580, 24'd7826962, 24'd8087494, 24'd8407614, 24'd8723974, 24'd8973965, 24'd9108115, 24'd9099876, 24'd8950878, 24'd8690607, 24'd8370572, 24'd8054106, 24'd7803837, 24'd7669293, 24'd7677100, 24'd7825713, 24'd8085722, 24'd8405671, 24'd8722244, 24'd8972790, 24'd9107728, 24'd9100353, 24'd8952125, 24'd8692378, 24'd8372515, 
24'd8055837, 24'd7805014, 24'd7669682, 24'd7676625, 24'd7824468, 24'd8083953, 24'd8403728, 24'd8720512, 24'd8971612, 24'd9107336, 24'd9100826, 24'd8953368, 24'd8694146, 24'd8374458, 24'd8057570, 24'd7806194, 24'd7670077, 24'd7676155, 24'd7823226, 24'd8082186, 24'd8401785, 24'd8718777, 24'd8970429, 24'd9106939, 24'd9101293, 24'd8954608, 24'd8695912, 24'd8376402, 24'd8059306, 24'd7807379, 
24'd7670476, 24'd7675690, 24'd7821989, 24'd8080421, 24'd8399842, 24'd8717040, 24'd8969242, 24'd9106537, 24'd9101756, 24'd8955843, 24'd8697676, 24'd8378345, 24'd8061044, 24'd7808568, 24'd7670881, 24'd7675230, 24'd7820755, 24'd8078658, 24'd8397898, 24'd8715301, 24'd8968051, 24'd9106130, 24'd9102213, 24'd8957075, 24'd8699438, 24'd8380288, 24'd8062785, 24'd7809761, 24'd7671290, 24'd7674775, 
24'd7819526, 24'd8076897, 24'd8395955, 24'd8713559, 24'd8966856, 24'd9105718, 24'd9102666, 24'd8958302, 24'd8701198, 24'd8382232, 24'd8064528, 24'd7810958, 24'd7671705, 24'd7674325, 24'd7818300, 24'd8075138, 24'd8394011, 24'd8711815, 24'd8965657, 24'd9105301, 24'd9103113, 24'd8959526, 24'd8702955, 24'd8384175, 24'd8066273, 24'd7812160, 24'd7672124, 24'd7673880, 24'd7817079, 24'd8073382, 
24'd8392068, 24'd8710069, 24'd8964453, 24'd9104879, 24'd9103556, 24'd8960745, 24'd8704710, 24'd8386119, 24'd8068020, 24'd7813365, 24'd7672549, 24'd7673440, 24'd7815861, 24'd8071628, 24'd8390124, 24'd8708321, 24'd8963246, 24'd9104452, 24'd9103993, 24'd8961961, 24'd8706463, 24'd8388062, 24'd8069769, 24'd7814574, 24'd7672979, 24'd7673005, 24'd7814648, 24'd8069876, 24'd8388181, 24'd8706570, 
24'd8962035, 24'd9104020, 24'd9104426, 24'd8963172, 24'd8708214, 24'd8390006, 24'd8071521, 24'd7815787, 24'd7673413, 24'd7672575, 24'd7813438, 24'd8068126, 24'd8386237, 24'd8704817, 24'd8960820, 24'd9103582, 24'd9104853, 24'd8964380, 24'd8709963, 24'd8391950, 24'd8073275, 24'd7817005, 24'd7673853, 24'd7672150, 24'd7812233, 24'd8066379, 24'd8384294, 24'd8703062, 24'd8959600, 24'd9103140, 
24'd9105275, 24'd8965583, 24'd8711709, 24'd8393893, 24'd8075031, 24'd7818226, 24'd7674298, 24'd7671730, 24'd7811031, 24'd8064634, 24'd8382350, 24'd8701305, 24'd8958377, 24'd9102693, 24'd9105693, 24'd8966783, 24'd8713453, 24'd8395837, 24'd8076790, 24'd7819451, 24'd7674747, 24'd7671315, 24'd7809834, 24'd8062891, 24'd8380407, 24'd8699545, 24'd8957150, 24'd9102241, 24'd9106105, 24'd8967978, 
24'd8715195, 24'd8397780, 24'd8078550, 24'd7820680, 24'd7675202, 24'd7670905, 24'd7808641, 24'd8061150, 24'd8378463, 24'd8697784, 24'd8955919, 24'd9101784, 24'd9106513, 24'd8969169, 24'd8716934, 24'd8399723, 24'd8080313, 24'd7821914, 24'd7675662, 24'd7670501, 24'd7807452, 24'd8059412, 24'd8376520, 24'd8696020, 24'd8954683, 24'd9101321, 24'd9106915, 24'd8970357, 24'd8718671, 24'd8401667, 
24'd8082078, 24'd7823151, 24'd7676127, 24'd7670101, 24'd7806266, 24'd8057676, 24'd8374577, 24'd8694254, 24'd8953444, 24'd9100854, 24'd9107312, 24'd8971540, 24'd8720406, 24'd8403610, 24'd8083845, 24'd7824392, 24'd7676596, 24'd7669706, 24'd7805085, 24'd8055942, 24'd8372633, 24'd8692486, 24'd8952201, 24'd9100382, 24'd9107704, 24'd8972719, 24'd8722138, 24'd8405553, 24'd8085614, 24'd7825637, 
24'd7677071, 24'd7669316, 24'd7803908, 24'd8054211, 24'd8370690, 24'd8690715, 24'd8950954, 24'd9099905, 24'd9108092, 24'd8973894, 24'd8723869, 24'd8407496, 24'd8087386, 24'd7826886, 24'd7677551, 24'd7668932, 24'd7802735, 24'd8052482, 24'd8368747, 24'd8688943, 24'd8949703, 24'd9099423, 24'd9108474, 24'd8975064, 24'd8725596, 24'd8409439, 24'd8089159, 24'd7828139, 24'd7678035, 24'd7668552, 
24'd7801567, 24'd8050756, 24'd8366805, 24'd8687169, 24'd8948448, 24'd9098936, 24'd9108851, 24'd8976231, 24'd8727322, 24'd8411382, 24'd8090935, 24'd7829396, 24'd7678525, 24'd7668178, 24'd7800402, 24'd8049031, 24'd8364862, 24'd8685392, 24'd8947189, 24'd9098443, 24'd9109223, 24'd8977394, 24'd8729045, 24'd8413324, 24'd8092712, 24'd7830657, 24'd7679020, 24'd7667808, 24'd7799241, 24'd8047309, 
24'd8362920, 24'd8683613, 24'd8945926, 24'd9097946, 24'd9109590, 24'd8978552, 24'd8730766, 24'd8415267, 24'd8094492, 24'd7831922, 24'd7679519, 24'd7667444, 24'd7798085, 24'd8045590, 24'd8360977, 24'd8681833, 24'd8944659, 24'd9097444, 24'd9109952, 24'd8979707, 24'd8732484, 24'd8417209, 24'd8096274, 24'd7833191, 24'd7680024, 24'd7667084, 24'd7796933, 24'd8043873, 24'd8359035, 24'd8680050, 
24'd8943389, 24'd9096937, 24'd9110309, 24'd8980857, 24'd8734200, 24'd8419151, 24'd8098057, 24'd7834463, 24'd7680533, 24'd7666730, 24'd7795785, 24'd8042158, 24'd8357093, 24'd8678265, 24'd8942114, 24'd9096425, 24'd9110660, 24'd8982003, 24'd8735913, 24'd8421093, 24'd8099843, 24'd7835740, 24'd7681048, 24'd7666381, 24'd7794641, 24'd8040446, 24'd8355152, 24'd8676478, 24'd8940836, 24'd9095908, 
24'd9111007, 24'd8983145, 24'd8737624, 24'd8423034, 24'd8101631, 24'd7837020, 24'd7681567, 24'd7666036, 24'd7793501, 24'd8038736, 24'd8353210, 24'd8674689, 24'd8939553, 24'd9095386, 24'd9111349, 24'd8984282, 24'd8739333, 24'd8424976, 24'd8103421, 24'd7838304, 24'd7682092, 24'd7665697, 24'd7792365, 24'd8037029, 24'd8351269, 24'd8672898, 24'd8938267, 24'd9094859, 24'd9111685, 24'd8985416, 
24'd8741039, 24'd8426917, 24'd8105213, 24'd7839592, 24'd7682621, 24'd7665363, 24'd7791234, 24'd8035324, 24'd8349328, 24'd8671105, 24'd8936977, 24'd9094327, 24'd9112017, 24'd8986545, 24'd8742743, 24'd8428857, 24'd8107007, 24'd7840884, 24'd7683155, 24'd7665034, 24'd7790107, 24'd8033621, 24'd8347387, 24'd8669311, 24'd8935683, 24'd9093791, 24'd9112344, 24'd8987670, 24'd8744444, 24'd8430798, 
24'd8108803, 24'd7842180, 24'd7683695, 24'd7664710, 24'd7788984, 24'd8031922, 24'd8345447, 24'd8667514, 24'd8934386, 24'd9093249, 24'd9112665, 24'd8988791, 24'd8746142, 24'd8432738, 24'd8110600, 24'd7843480, 24'd7684239, 24'd7664391, 24'd7787865, 24'd8030224, 24'd8343507, 24'd8665715, 24'd8933084, 24'd9092702, 24'd9112981, 24'd8989908, 24'd8747839, 24'd8434678, 24'd8112400, 24'd7844783, 
24'd7684788, 24'd7664077, 24'd7786750, 24'd8028529, 24'd8341567, 24'd8663914, 24'd8931779, 24'd9092151, 24'd9113293, 24'd8991021, 24'd8749532, 24'd8436618, 24'd8114202, 24'd7846090, 24'd7685342, 24'd7663769, 24'd7785640, 24'd8026837, 24'd8339628, 24'd8662112, 24'd8930470, 24'd9091594, 24'd9113599, 24'd8992129, 24'd8751223, 24'd8438557, 24'd8116005, 24'd7847401, 24'd7685901, 24'd7663465, 
24'd7784534, 24'd8025147, 24'd8337689, 24'd8660307, 24'd8929157, 24'd9091033, 24'd9113900, 24'd8993233, 24'd8752912, 24'd8440496, 24'd8117811, 24'd7848716, 24'd7686465, 24'd7663167, 24'd7783432, 24'd8023460, 24'd8335750, 24'd8658501, 24'd8927840, 24'd9090466, 24'd9114196, 24'd8994333, 24'd8754598, 24'd8442434, 24'd8119618, 24'd7850035, 24'd7687034, 24'd7662873, 24'd7782334, 24'd8021775, 
24'd8333812, 24'd8656692, 24'd8926519, 24'd9089895, 24'd9114487, 24'd8995428, 24'd8756281, 24'd8444372, 24'd8121428, 24'd7851357, 24'd7687608, 24'd7662585, 24'd7781240, 24'd8020093, 24'd8331874, 24'd8654882, 24'd8925195, 24'd9089319, 24'd9114773, 24'd8996520, 24'd8757962, 24'd8446310, 24'd8123239, 24'd7852683, 24'd7688186, 24'd7662301, 24'd7780151, 24'd8018413, 24'd8329936, 24'd8653070, 
24'd8923867, 24'd9088737, 24'd9115053, 24'd8997607, 24'd8759641, 24'd8448248, 24'd8125052, 24'd7854013, 24'd7688770, 24'd7662023, 24'd7779066, 24'd8016736, 24'd8327999, 24'd8651256, 24'd8922535, 24'd9088151, 24'd9115329, 24'd8998690, 24'd8761316, 24'd8450184, 24'd8126867, 24'd7855347, 24'd7689359, 24'd7661750, 24'd7777986, 24'd8015062, 24'd8326062, 24'd8649440, 24'd8921200, 24'd9087560, 
24'd9115599, 24'd8999768, 24'd8762989, 24'd8452121, 24'd8128683, 24'd7856684, 24'd7689952, 24'd7661482, 24'd7776909, 24'd8013390, 24'd8324126, 24'd8647623, 24'd8919860, 24'd9086964, 24'd9115865, 24'd9000842, 24'd8764660, 24'd8454057, 24'd8130502, 24'd7858026, 24'd7690550, 24'd7661219, 24'd7775837, 24'd8011721, 24'd8322190, 24'd8645803, 24'd8918517, 24'd9086364, 24'd9116125, 24'd9001912, 
24'd8766328, 24'd8455993, 24'd8132322, 24'd7859370, 24'd7691154, 24'd7660962, 24'd7774769, 24'd8010055, 24'd8320255, 24'd8643982, 24'd8917171, 24'd9085758, 24'd9116380, 24'd9002978, 24'd8767993, 24'd8457928, 24'd8134144, 24'd7860719, 24'd7691762, 24'd7660709, 24'd7773706, 24'd8008391, 24'd8318320, 24'd8642159, 24'd8915820, 24'd9085147, 24'd9116631, 24'd9004039, 24'd8769655, 24'd8459862, 
24'd8135968, 24'd7862071, 24'd7692375, 24'd7660461, 24'd7772647, 24'd8006730, 24'd8316385, 24'd8640334, 24'd8914466, 24'd9084532, 24'd9116876, 24'd9005096, 24'd8771315, 24'd8461797, 24'd8137794, 24'd7863427, 24'd7692993, 24'd7660219, 24'd7771592, 24'd8005071, 24'd8314452, 24'd8638507, 24'd8913108, 24'd9083912, 24'd9117116, 24'd9006149, 24'd8772972, 24'd8463730, 24'd8139622, 24'd7864787, 
24'd7693615, 24'd7659981, 24'd7770541, 24'd8003415, 24'd8312518, 24'd8636679, 24'd8911747, 24'd9083287, 24'd9117350, 24'd9007197, 24'd8774627, 24'd8465663, 24'd8141451, 24'd7866150, 24'd7694243, 24'd7659749, 24'd7769495, 24'd8001762, 24'd8310585, 24'd8634849, 24'd8910382, 24'd9082656, 24'd9117580, 24'd9008241, 24'd8776278, 24'd8467596, 24'd8143282, 24'd7867517, 24'd7694875, 24'd7659522, 
24'd7768453, 24'd8000112, 24'd8308653, 24'd8633017, 24'd8909013, 24'd9082022, 24'd9117805, 24'd9009281, 24'd8777927, 24'd8469528, 24'd8145114, 24'd7868888, 24'd7695513, 24'd7659300, 24'd7767416, 24'd7998464, 24'd8306721, 24'd8631184, 24'd8907641, 24'd9081382, 24'd9118024, 24'd9010316, 24'd8779574, 24'd8471459, 24'd8146949, 24'd7870262, 24'd7696155, 24'd7659083, 24'd7766383, 24'd7996819, 
24'd8304790, 24'd8629348, 24'd8906264, 24'd9080737, 24'd9118239, 24'd9011347, 24'd8781217, 24'd8473390, 24'd8148785, 24'd7871640, 24'd7696802, 24'd7658871, 24'd7765354, 24'd7995177, 24'd8302860, 24'd8627511, 24'd8904885, 24'd9080088, 24'd9118448, 24'd9012374, 24'd8782858, 24'd8475320, 24'd8150623, 24'd7873022, 24'd7697454, 24'd7658664, 24'd7764329, 24'd7993538, 24'd8300930, 24'd8625673, 
24'd8903501, 24'd9079433, 24'd9118652, 24'd9013396, 24'd8784496, 24'd8477250, 24'd8152462, 24'd7874407, 24'd7698111, 24'd7658463, 24'd7763309, 24'd7991901, 24'd8299000, 24'd8623833, 24'd8902114, 24'd9078774, 24'd9118851, 24'd9014414, 24'd8786131, 24'd8479179, 24'd8154303, 24'd7875795, 24'd7698772, 24'd7658266, 24'd7762294, 24'd7990267, 24'd8297072, 24'd8621991, 24'd8900724, 24'd9078110, 
24'd9119045, 24'd9015428, 24'd8787764, 24'd8481108, 24'd8156146, 24'd7877188, 24'd7699439, 24'd7658075, 24'd7761282, 24'd7988636, 24'd8295143, 24'd8620147, 24'd8899330, 24'd9077441, 24'd9119234, 24'd9016437, 24'd8789393, 24'd8483035, 24'd8157990, 24'd7878584, 24'd7700110, 24'd7657889, 24'd7760275, 24'd7987008, 24'd8293216, 24'd8618302, 24'd8897932, 24'd9076767, 24'd9119417, 24'd9017441, 
24'd8791020, 24'd8484962, 24'd8159836, 24'd7879983, 24'd7700786, 24'd7657708, 24'd7759273, 24'd7985382, 24'd8291289, 24'd8616455, 24'd8896531, 24'd9076089, 24'd9119596, 24'd9018442, 24'd8792644, 24'd8486889, 24'd8161684, 24'd7881386, 24'd7701467, 24'd7657532, 24'd7758275, 24'd7983760, 24'd8289363, 24'd8614607, 24'd8895126, 24'd9075406, 24'd9119769, 24'd9019437, 24'd8794265, 24'd8488815, 
24'd8163533, 24'd7882793, 24'd7702153, 24'd7657361, 24'd7757281, 24'd7982140, 24'd8287438, 24'd8612757, 24'd8893717, 24'd9074717, 24'd9119938, 24'd9020429, 24'd8795884, 24'd8490740, 24'd8165384, 24'd7884203, 24'd7702843, 24'd7657195, 24'd7756292, 24'd7980523, 24'd8285513, 24'd8610905, 24'd8892305, 24'd9074024, 24'd9120101, 24'd9021416, 24'd8797499, 24'd8492664, 24'd8167236, 24'd7885617, 
24'd7703539, 24'd7657035, 24'd7755307, 24'd7978909, 24'd8283589, 24'd8609052, 24'd8890890, 24'd9073327, 24'd9120259, 24'd9022398, 24'd8799112, 24'd8494587, 24'd8169090, 24'd7887034, 24'd7704239, 24'd7656879, 24'd7754327, 24'd7977298, 24'd8281666, 24'd8607198, 24'd8889471, 24'd9072624, 24'd9120412, 24'd9023377, 24'd8800722, 24'd8496510, 24'd8170945, 24'd7888455, 24'd7704944, 24'd7656729, 
24'd7753351, 24'd7975689, 24'd8279744, 24'd8605342, 24'd8888048, 24'd9071917, 24'd9120559, 24'd9024350, 24'd8802329, 24'd8498432, 24'd8172802, 24'd7889879, 24'd7705654, 24'd7656584, 24'd7752380, 24'd7974084, 24'd8277822, 24'd8603484, 24'd8886622, 24'd9071205, 24'd9120702, 24'd9025319, 24'd8803933, 24'd8500354, 24'd8174660, 24'd7891307, 24'd7706368, 24'd7656444, 24'd7751413, 24'd7972482, 
24'd8275901, 24'd8601625, 24'd8885193, 24'd9070488, 24'd9120840, 24'd9026284, 24'd8805534, 24'd8502274, 24'd8176520, 24'd7892738, 24'd7707088, 24'd7656309, 24'd7750450, 24'd7970882, 24'd8273981, 24'd8599764, 24'd8883760, 24'd9069766, 24'd9120972, 24'd9027244, 24'd8807132, 24'd8504194, 24'd8178382, 24'd7894173, 24'd7707812, 24'd7656179, 24'd7749492, 24'd7969285, 24'd8272061, 24'd8597902, 
24'd8882323, 24'd9069039, 24'd9121099, 24'd9028200, 24'd8808727, 24'd8506113, 24'd8180245, 24'd7895611, 24'd7708541, 24'd7656054, 24'd7748539, 24'd7967692, 24'd8270143, 24'd8596038, 24'd8880884, 24'd9068308, 24'd9121221, 24'd9029152, 24'd8810319, 24'd8508031, 24'd8182109, 24'd7897053, 24'd7709274, 24'd7655935, 24'd7747590, 24'd7966101, 24'd8268225, 24'd8594173, 24'd8879440, 24'd9067572, 
24'd9121338, 24'd9030098, 24'd8811909, 24'd8509948, 24'd8183975, 24'd7898498, 24'd7710013, 24'd7655820, 24'd7746645, 24'd7964513, 24'd8266308, 24'd8592307, 24'd8877993, 24'd9066831, 24'd9121450, 24'd9031041, 24'd8813495, 24'd8511865, 24'd8185842, 24'd7899946, 24'd7710756, 24'd7655711, 24'd7745705, 24'd7962928, 24'd8264392, 24'd8590439, 24'd8876543, 24'd9066086, 24'd9121557, 24'd9031978, 
24'd8815078, 24'd8513780, 24'd8187711, 24'd7901398, 24'd7711504, 24'd7655607, 24'd7744769, 24'd7961346, 24'd8262477, 24'd8588569, 24'd8875089, 24'd9065335, 24'd9121658, 24'd9032912, 24'd8816659, 24'd8515695, 24'd8189581, 24'd7902854, 24'd7712256, 24'd7655508, 24'd7743838, 24'd7959767, 24'd8260563, 24'd8586699, 24'd8873632, 24'd9064580, 24'd9121755, 24'd9033841, 24'd8818236, 24'd8517609, 
24'd8191452, 24'd7904313, 24'd7713014, 24'd7655414, 24'd7742912, 24'd7958192, 24'd8258650, 24'd8584827, 24'd8872172, 24'd9063821, 24'd9121846, 24'd9034765, 24'd8819810, 24'd8519521, 24'd8193325, 24'd7905775, 24'd7713776, 24'd7655325, 24'd7741990, 24'd7956619, 24'd8256737, 24'd8582953, 24'd8870708, 24'd9063056, 24'd9121932, 24'd9035685, 24'd8821382, 24'd8521433, 24'd8195199, 24'd7907240, 
24'd7714543, 24'd7655242, 24'd7741072, 24'd7955049, 24'd8254826, 24'd8581078, 24'd8869241, 24'd9062287, 24'd9122013, 24'd9036600, 24'd8822950, 24'd8523344, 24'd8197075, 24'd7908709, 24'd7715315, 24'd7655163, 24'd7740159, 24'd7953482, 24'd8252915, 24'd8579202, 24'd8867770, 24'd9061513, 24'd9122089, 24'd9037510, 24'd8824515, 24'd8525255, 24'd8198952, 24'd7910182, 24'd7716091, 24'd7655090, 
24'd7739251, 24'd7951918, 24'd8251006, 24'd8577324, 24'd8866296, 24'd9060734, 24'd9122160, 24'd9038416, 24'd8826077, 24'd8527164, 24'd8200830, 24'd7911657, 24'd7716872, 24'd7655022, 24'd7738347, 24'd7950358, 24'd8249097, 24'd8575445, 24'd8864819, 24'd9059951, 24'd9122225, 24'd9039318, 24'd8827636, 24'd8529072, 24'd8202710, 24'd7913136, 24'd7717658, 24'd7654959, 24'd7737448, 24'd7948800, 
24'd8247189, 24'd8573565, 24'd8863338, 24'd9059163, 24'd9122286, 24'd9040215, 24'd8829192, 24'd8530979, 24'd8204590, 24'd7914619, 24'd7718448, 24'd7654901, 24'd7736553, 24'd7947246, 24'd8245283, 24'd8571684, 24'd8861854, 24'd9058370, 24'd9122341, 24'd9041107, 24'd8830745, 24'd8532885, 24'd8206473, 24'd7916104, 24'd7719243, 24'd7654848, 24'd7735663, 24'd7945694, 24'd8243377, 24'd8569801, 
24'd8860367, 24'd9057572, 24'd9122391, 24'd9041995, 24'd8832295, 24'd8534790, 24'd8208356, 24'd7917593, 24'd7720043, 24'd7654801, 24'd7734778, 24'd7944146, 24'd8241473, 24'd8567917, 24'd8858876, 24'd9056770, 24'd9122436, 24'd9042879, 24'd8833842, 24'd8536694, 24'd8210241, 24'd7919085, 24'd7720848, 24'd7654758, 24'd7733897, 24'd7942601, 24'd8239569, 24'd8566031, 24'd8857382, 24'd9055963, 
24'd9122476, 24'd9043757, 24'd8835386, 24'd8538598, 24'd8212127, 24'd7920581, 24'd7721657, 24'd7654721, 24'd7733020, 24'd7941059, 24'd8237666, 24'd8564145, 24'd8855885, 24'd9055152, 24'd9122510, 24'd9044631, 24'd8836926, 24'd8540500, 24'd8214014, 24'd7922080, 24'd7722471, 24'd7654689, 24'd7732148, 24'd7939520, 24'd8235765, 24'd8562257, 24'd8854384, 24'd9054335, 24'd9122540, 24'd9045501, 
24'd8838463, 24'd8542401, 24'd8215902, 24'd7923582, 24'd7723289, 24'd7654662, 24'd7731281, 24'd7937984, 24'd8233864, 24'd8560368, 24'd8852881, 24'd9053515, 24'd9122564, 24'd9046366, 24'd8839998, 24'd8544300, 24'd8217792, 24'd7925087, 24'd7724113, 24'd7654640, 24'd7730419, 24'd7936451, 24'd8231965, 24'd8558478, 24'd8851374, 24'd9052689, 24'd9122584, 24'd9047226, 24'd8841529, 24'd8546199, 
24'd8219683, 24'd7926596, 24'd7724941, 24'd7654624, 24'd7729561, 24'd7934922, 24'd8230067, 24'd8556586, 24'd8849863, 24'd9051859, 24'd9122598, 24'd9048082, 24'd8843057, 24'd8548097, 24'd8221575, 24'd7928108, 24'd7725773, 24'd7654612, 24'd7728707, 24'd7933396, 24'd8228170, 24'd8554694, 24'd8848350, 24'd9051024, 24'd9122607, 24'd9048933, 24'd8844581, 24'd8549994, 24'd8223468, 24'd7929623, 
24'd7726610, 24'd7654606, 24'd7727859, 24'd7931873, 24'd8226274, 24'd8552800, 24'd8846833, 24'd9050184, 24'd9122611, 24'd9049779, 24'd8846103, 24'd8551889, 24'd8225362, 24'd7931141, 24'd7727452, 24'd7654604, 24'd7727015, 24'd7930353, 24'd8224379, 24'd8550905, 24'd8845313, 24'd9049340, 24'd9122609, 24'd9050621, 24'd8847621, 24'd8553783, 24'd8227258, 24'd7932663, 24'd7728299, 24'd7654608, 
24'd7726175, 24'd7928836, 24'd8222485, 24'd8549009, 24'd8843790, 24'd9048491, 24'd9122603, 24'd9051458, 24'd8849136, 24'd8555676, 24'd8229154, 24'd7934188, 24'd7729150, 24'd7654617, 24'd7725340, 24'd7927323, 24'd8220592, 24'd8547112, 24'd8842264, 24'd9047638, 24'd9122591, 24'd9052290, 24'd8850648, 24'd8557568, 24'd8231052, 24'd7935715, 24'd7730005, 24'd7654632, 24'd7724510, 24'd7925813, 
24'd8218701, 24'd8545214, 24'd8840734, 24'd9046780, 24'd9122574, 24'd9053118, 24'd8852156, 24'd8559459, 24'd8232951, 24'd7937247, 24'd7730866, 24'd7654651, 24'd7723685, 24'd7924306, 24'd8216811, 24'd8543314, 24'd8839202, 24'd9045917, 24'd9122552, 24'd9053941, 24'd8853662, 24'd8561349, 24'd8234851, 24'd7938781, 24'd7731731, 24'd7654675, 24'd7722864, 24'd7922802, 24'd8214922, 24'd8541414, 
24'd8837666, 24'd9045050, 24'd9122525, 24'd9054760, 24'd8855164, 24'd8563237, 24'd8236752, 24'd7940318, 24'd7732600, 24'd7654705, 24'd7722048, 24'd7921301, 24'd8213034, 24'd8539512, 24'd8836127, 24'd9044178, 24'd9122493, 24'd9055573, 24'd8856663, 24'd8565124, 24'd8238654, 24'd7941859, 24'd7733475, 24'd7654740, 24'd7721236, 24'd7919804, 24'd8211148, 24'd8537610, 24'd8834585, 24'd9043302, 
24'd9122456, 24'd9056383, 24'd8858158, 24'd8567010, 24'd8240557, 24'd7943402, 24'd7734353, 24'd7654780, 24'd7720430, 24'd7918310, 24'd8209262, 24'd8535706, 24'd8833040, 24'd9042421, 24'd9122413, 24'd9057187, 24'd8859650, 24'd8568895, 24'd8242461, 24'd7944949, 24'd7735237, 24'd7654825, 24'd7719627, 24'd7916820, 24'd8207378, 24'd8533802, 24'd8831491, 24'd9041535, 24'd9122366, 24'd9057987, 
24'd8861139, 24'd8570778, 24'd8244366, 24'd7946499, 24'd7736125, 24'd7654875, 24'd7718830, 24'd7915333, 24'd8205495, 24'd8531896, 24'd8829940, 24'd9040645, 24'd9122313, 24'd9058782, 24'd8862625, 24'd8572660, 24'd8246272, 24'd7948052, 24'd7737017, 24'd7654930, 24'd7718037, 24'd7913849, 24'd8203614, 24'd8529989, 24'd8828385, 24'd9039750, 24'd9122255, 24'd9059572, 24'd8864107, 24'd8574541, 
24'd8248180, 24'd7949608, 24'd7737914, 24'd7654991, 24'd7717249, 24'd7912368, 24'd8201734, 24'd8528082, 24'd8826828, 24'd9038851, 24'd9122192, 24'd9060358, 24'd8865586, 24'd8576421, 24'd8250088, 24'd7951167, 24'd7738816, 24'd7655057, 24'd7716466, 24'd7910891, 24'd8199855, 24'd8526173, 24'd8825267, 24'd9037947, 24'd9122124, 24'd9061139, 24'd8867062, 24'd8578299, 24'd8251997, 24'd7952730, 
24'd7739722, 24'd7655127, 24'd7715687, 24'd7909417, 24'd8197977, 24'd8524263, 24'd8823703, 24'd9037038, 24'd9122050, 24'd9061915, 24'd8868534, 24'd8580176, 24'd8253907, 24'd7954295, 24'd7740633, 24'd7655203, 24'd7714913, 24'd7907946, 24'd8196101, 24'd8522353, 24'd8822136, 24'd9036125, 24'd9121972, 24'd9062687, 24'd8870003, 24'd8582051, 24'd8255818, 24'd7955863, 24'd7741548, 24'd7655284, 
24'd7714144, 24'd7906479, 24'd8194226, 24'd8520441, 24'd8820566, 24'd9035208, 24'd9121888, 24'd9063454, 24'd8871468, 24'd8583926, 24'd8257730, 24'd7957435, 24'd7742468, 24'd7655371, 24'd7713380, 24'd7905015, 24'd8192353, 24'd8518529, 24'd8818993, 24'd9034286, 24'd9121799, 24'd9064216, 24'd8872930, 24'd8585798, 24'd8259643, 24'd7959009, 24'd7743392, 24'd7655462, 24'd7712620, 24'd7903555, 
24'd8190481, 24'd8516615, 24'd8817418, 24'd9033359, 24'd9121705, 24'd9064973, 24'd8874389, 24'd8587670, 24'd8261557, 24'd7960587, 24'd7744321, 24'd7655559, 24'd7711865, 24'd7902098, 24'd8188610, 24'd8514701, 24'd8815839, 24'd9032428, 24'd9121606, 24'd9065725, 24'd8875844, 24'd8589540, 24'd8263471, 24'd7962167, 24'd7745254, 24'd7655660, 24'd7711115, 24'd7900644, 24'd8186741, 24'd8512786, 
24'd8814257, 24'd9031492, 24'd9121502, 24'd9066473, 24'd8877296, 24'd8591409, 24'd8265387, 24'd7963750, 24'd7746192, 24'd7655767, 24'd7710370, 24'd7899194, 24'd8184873, 24'd8510870, 24'd8812672, 24'd9030552, 24'd9121393, 24'd9067216, 24'd8878745, 24'd8593276, 24'd8267303, 24'd7965337, 24'd7747135, 24'd7655879, 24'd7709629, 24'd7897747, 24'd8183006, 24'd8508953, 24'd8811084, 24'd9029607, 
24'd9121278, 24'd9067955, 24'd8880190, 24'd8595141, 24'd8269221, 24'd7966926, 24'd7748082, 24'd7655996, 24'd7708893, 24'd7896304, 24'd8181141, 24'd8507035, 24'd8809493, 24'd9028658, 24'd9121159, 24'd9068688, 24'd8881631, 24'd8597006, 24'd8271139, 24'd7968518, 24'd7749033, 24'd7656118, 24'd7708162, 24'd7894864, 24'd8179278, 24'd8505117, 24'd8807899, 24'd9027705, 24'd9121034, 24'd9069417, 
24'd8883069, 24'd8598869, 24'd8273058, 24'd7970114, 24'd7749989, 24'd7656246, 24'd7707435, 24'd7893428, 24'd8177415, 24'd8503198, 24'd8806303, 24'd9026747, 24'd9120904, 24'd9070141, 24'd8884504, 24'd8600730, 24'd8274977, 24'd7971712, 24'd7750949, 24'd7656378, 24'd7706714, 24'd7891995, 24'd8175555, 24'd8501277, 24'd8804703, 24'd9025784, 24'd9120769, 24'd9070860, 24'd8885935, 24'd8602590, 
24'd8276898, 24'd7973313, 24'd7751914, 24'd7656516, 24'd7705997, 24'd7890565, 24'd8173696, 24'd8499357, 24'd8803100, 24'd9024817, 24'd9120629, 24'd9071575, 24'd8887363, 24'd8604448, 24'd8278819, 24'd7974917, 24'd7752883, 24'd7656658, 24'd7705285, 24'd7889139, 24'd8171838, 24'd8497435, 24'd8801495, 24'd9023845, 24'd9120483, 24'd9072285, 24'd8888787, 24'd8606305, 24'd8280741, 24'd7976524, 
24'd7753857, 24'd7656806, 24'd7704577, 24'd7887717, 24'd8169982, 24'd8495512, 24'd8799887, 24'd9022869, 24'd9120333, 24'd9072989, 24'd8890208, 24'd8608161, 24'd8282664, 24'd7978134, 24'd7754835, 24'd7656959, 24'd7703875, 24'd7886298, 24'd8168127, 24'd8493589, 24'd8798275, 24'd9021889, 24'd9120177, 24'd9073689, 24'd8891625, 24'd8610014, 24'd8284588, 24'd7979746, 24'd7755818, 24'd7657117, 
24'd7703177, 24'd7884883, 24'd8166274, 24'd8491665, 24'd8796661, 24'd9020904, 24'd9120017, 24'd9074385, 24'd8893039, 24'd8611867, 24'd8286512, 24'd7981362, 24'd7756805, 24'd7657281, 24'd7702484, 24'd7883471, 24'd8164423, 24'd8489740, 24'd8795044, 24'd9019915, 24'd9119851, 24'd9075075, 24'd8894449, 24'd8613717, 24'd8288437, 24'd7982980, 24'd7757796, 24'd7657449, 24'd7701796, 24'd7882062, 
24'd8162573, 24'd8487815, 24'd8793424, 24'd9018921, 24'd9119680, 24'd9075761, 24'd8895855, 24'd8615567, 24'd8290363, 24'd7984602, 24'd7758792, 24'd7657622, 24'd7701113, 24'd7880658, 24'd8160724, 24'd8485889, 24'd8791802, 24'd9017923, 24'd9119504, 24'd9076442, 24'd8897258, 24'd8617414, 24'd8292289, 24'd7986226, 24'd7759793, 24'd7657801, 24'd7700435, 24'd7879256, 24'd8158878, 24'd8483962, 
24'd8790176, 24'd9016920, 24'd9119323, 24'd9077118, 24'd8898658, 24'd8619260, 24'd8294216, 24'd7987853, 24'd7760798, 24'd7657985, 24'd7699761, 24'd7877859, 24'd8157033, 24'd8482035, 24'd8788548, 24'd9015913, 24'd9119136, 24'd9077789, 24'd8900054, 24'd8621104, 24'd8296144, 24'd7989482, 24'd7761807, 24'd7658174, 24'd7699092, 24'd7876465, 24'd8155189, 24'd8480107, 24'd8786917, 24'd9014902, 
24'd9118945, 24'd9078455, 24'd8901446, 24'd8622947, 24'd8298073, 24'd7991115, 24'd7762820, 24'd7658368, 24'd7698428, 24'd7875074, 24'd8153347, 24'd8478178, 24'd8785283, 24'd9013886, 24'd9118748, 24'd9079117, 24'd8902835, 24'd8624788, 24'd8300002, 24'd7992750, 24'd7763838, 24'd7658567, 24'd7697769, 24'd7873687, 24'd8151507, 24'd8476249, 24'd8783646, 24'd9012866, 24'd9118547, 24'd9079773, 
24'd8904220, 24'd8626627, 24'd8301931, 24'd7994388, 24'd7764860, 24'd7658771, 24'd7697115, 24'd7872304, 24'd8149669, 24'd8474319, 24'd8782007, 24'd9011842, 24'd9118340, 24'd9080425, 24'd8905601, 24'd8628465, 24'd8303862, 24'd7996029, 24'd7765887, 24'd7658980, 24'd7696466, 24'd7870924, 24'd8147832, 24'd8472388, 24'd8780364, 24'd9010813, 24'd9118128, 24'd9081072, 24'd8906979, 24'd8630301, 
24'd8305792, 24'd7997673, 24'd7766918, 24'd7659195, 24'd7695821, 24'd7869548, 24'd8145996, 24'd8470457, 24'd8778719, 24'd9009780, 24'd9117911, 24'd9081714, 24'd8908353, 24'd8632136, 24'd8307724, 24'd7999319, 24'd7767954, 24'd7659415, 24'd7695181, 24'd7868176, 24'd8144163, 24'd8468525, 24'd8777072, 24'd9008742, 24'd9117689, 24'd9082352, 24'd8909724, 24'd8633968, 24'd8309656, 24'd8000968, 
24'd7768993, 24'd7659639, 24'd7694546, 24'd7866807, 24'd8142331, 24'd8466593, 24'd8775421, 24'd9007700, 24'd9117462, 24'd9082984, 24'd8911091, 24'd8635799, 24'd8311589, 24'd8002620, 24'd7770038, 24'd7659869, 24'd7693917, 24'd7865442, 24'd8140501, 24'd8464660, 24'd8773768, 24'd9006654, 24'd9117229, 24'd9083612, 24'd8912454, 24'd8637628, 24'd8313522, 24'd8004274, 24'd7771086, 24'd7660104, 
24'd7693291, 24'd7864081, 24'd8138673, 24'd8462727, 24'd8772112, 24'd9005603, 24'd9116992, 24'd9084234, 24'd8913814, 24'd8639456, 24'd8315455, 24'd8005932, 24'd7772139, 24'd7660344, 24'd7692671, 24'd7862723, 24'd8136846, 24'd8460793, 24'd8770454, 24'd9004548, 24'd9116749, 24'd9084852, 24'd8915170, 24'd8641281, 24'd8317389, 24'd8007591, 24'd7773196, 24'd7660589, 24'd7692056, 24'd7861369, 
24'd8135021, 24'd8458858, 24'd8768793, 24'd9003489, 24'd9116501, 24'd9085465, 24'd8916522, 24'd8643105, 24'd8319324, 24'd8009254, 24'd7774257, 24'd7660839, 24'd7691445, 24'd7860019, 24'd8133198, 24'd8456923, 24'd8767129, 24'd9002425, 24'd9116249, 24'd9086073, 24'd8917870, 24'd8644927, 24'd8321259, 24'd8010919, 24'd7775323, 24'd7661095, 24'd7690840, 24'd7858672, 24'd8131377, 24'd8454988, 
24'd8765462, 24'd9001358, 24'd9115991, 24'd9086676, 24'd8919215, 24'd8646748, 24'd8323195, 24'd8012587, 24'd7776393, 24'd7661355, 24'd7690239, 24'd7857329, 24'd8129558, 24'd8453052, 24'd8763793, 24'd9000285, 24'd9115728, 24'd9087274, 24'd8920556, 24'd8648566, 24'd8325131, 24'd8014258, 24'd7777467, 24'd7661621, 24'd7689643, 24'd7855990, 24'd8127740, 24'd8451116, 24'd8762121, 24'd8999209, 
24'd9115460, 24'd9087868, 24'd8921893, 24'd8650383, 24'd8327067, 24'd8015931, 24'd7778546, 24'd7661891, 24'd7689052, 24'd7854654, 24'd8125924, 24'd8449179, 24'd8760447, 24'd8998128, 24'd9115186, 24'd9088456, 24'd8923227, 24'd8652198, 24'd8329004, 24'd8017606, 24'd7779629, 24'd7662167, 24'd7688467, 24'd7853323, 24'd8124111, 24'd8447242, 24'd8758770, 24'd8997043, 24'd9114908, 24'd9089040, 
24'd8924557, 24'd8654011, 24'd8330942, 24'd8019285, 24'd7780716, 24'd7662448, 24'd7687885, 24'd7851995, 24'd8122298, 24'd8445304, 24'd8757090, 24'd8995954, 24'd9114625, 24'd9089618, 24'd8925883, 24'd8655822, 24'd8332880, 24'd8020966, 24'd7781807, 24'd7662734, 24'd7687309, 24'd7850670, 24'd8120488, 24'd8443366, 24'd8755408, 24'd8994860, 24'd9114336, 24'd9090192, 24'd8927205, 24'd8657631, 
24'd8334818, 24'd8022649, 24'd7782903, 24'd7663025, 24'd7686738, 24'd7849350, 24'd8118680, 24'd8441428, 24'd8753723, 24'd8993762, 24'd9114043, 24'd9090761, 24'd8928524, 24'd8659439, 24'd8336756, 24'd8024335, 24'd7784003, 24'd7663321, 24'd7686172, 24'd7848033, 24'd8116874, 24'd8439489, 24'd8752036, 24'd8992660, 24'd9113744, 24'd9091325, 24'd8929839, 24'd8661244, 24'd8338695, 24'd8026024, 
24'd7785107, 24'd7663622, 24'd7685610, 24'd7846720, 24'd8115069, 24'd8437550, 24'd8750346, 24'd8991554, 24'd9113440, 24'd9091884, 24'd8931150, 24'd8663048, 24'd8340634, 24'd8027715, 24'd7786216, 24'd7663928, 24'd7685054, 24'd7845411, 24'd8113266, 24'd8435611, 24'd8748654, 24'd8990444, 24'd9113132, 24'd9092438, 24'd8932457, 24'd8664849, 24'd8342574, 24'd8029409, 24'd7787328, 24'd7664240, 
24'd7684502, 24'd7844106, 24'd8111466, 24'd8433671, 24'd8746959, 24'd8989329, 24'd9112818, 24'd9092987, 24'd8933760, 24'd8666649, 24'd8344514, 24'd8031105, 24'd7788445, 24'd7664556, 24'd7683956, 24'd7842805, 24'd8109667, 24'd8431731, 24'd8745261, 24'd8988210, 24'd9112499, 24'd9093531, 24'd8935060, 24'd8668447, 24'd8346454, 24'd8032804, 24'd7789566, 24'd7664878, 24'd7683414, 24'd7841507, 
24'd8107870, 24'd8429791, 24'd8743561, 24'd8987087, 24'd9112175, 24'd9094070, 24'd8936355, 24'd8670242, 24'd8348395, 24'd8034505, 24'd7790691, 24'd7665204, 24'd7682877, 24'd7840213, 24'd8106075, 24'd8427850, 24'd8741859, 24'd8985960, 24'd9111846, 24'd9094604, 24'd8937647, 24'd8672036, 24'd8350335, 24'd8036208, 24'd7791821, 24'd7665536, 24'd7682346, 24'd7838923, 24'd8104283, 24'd8425909, 
24'd8740154, 24'd8984828, 24'd9111511, 24'd9095133, 24'd8938935, 24'd8673828, 24'd8352276, 24'd8037915, 24'd7792954, 24'd7665873, 24'd7681819, 24'd7837637, 24'd8102492, 24'd8423968, 24'd8738446, 24'd8983692, 24'd9111172, 24'd9095658, 24'd8940219, 24'd8675618, 24'd8354218, 24'd8039623, 24'd7794092, 24'd7666214, 24'd7681297, 24'd7836355, 24'd8100703, 24'd8422026, 24'd8736737, 24'd8982552, 
24'd9110828, 24'd9096177, 24'd8941500, 24'd8677406, 24'd8356159, 24'd8041334, 24'd7795234, 24'd7666561, 24'd7680780, 24'd7835077, 24'd8098916, 24'd8420085, 24'd8735024, 24'd8981408, 24'd9110478, 24'd9096691, 24'd8942776, 24'd8679192, 24'd8358101, 24'd8043048, 24'd7796380, 24'd7666913, 24'd7680268, 24'd7833802, 24'd8097131, 24'd8418143, 24'd8733310, 24'd8980260, 24'd9110124, 24'd9097201, 
24'd8944049, 24'd8680975, 24'd8360043, 24'd8044764, 24'd7797530, 24'd7667270, 24'd7679761, 24'd7832532, 24'd8095349, 24'd8416201, 24'd8731592, 24'd8979108, 24'd9109764, 24'd9097705, 24'd8945317, 24'd8682757, 24'd8361985, 24'd8046482, 24'd7798685, 24'd7667632, 24'd7679259, 24'd7831265, 24'd8093568, 24'd8414258, 24'd8729873, 24'd8977951, 24'd9109400, 24'd9098205, 24'd8946582, 24'd8684537, 
24'd8363928, 24'd8048203, 24'd7799843, 24'd7667999, 24'd7678762, 24'd7830002, 24'd8091789, 24'd8412316, 24'd8728151, 24'd8976791, 24'd9109030, 24'd9098699, 24'd8947843, 24'd8686314, 24'd8365870, 24'd8049926, 24'd7801006, 24'd7668371, 24'd7678270, 24'd7828743, 24'd8090013, 24'd8410373, 24'd8726427, 24'd8975626, 24'd9108656, 24'd9099189, 24'd8949100, 24'd8688090, 24'd8367813, 24'd8051651, 
24'd7802173, 24'd7668749, 24'd7677783, 24'd7827488, 24'd8088238, 24'd8408431, 24'd8724700, 24'd8974457, 24'd9108276, 24'd9099674, 24'd8950353, 24'd8689863, 24'd8369756, 24'd8053379, 24'd7803344, 24'd7669131, 24'd7677301, 24'd7826237, 24'd8086466, 24'd8406488, 24'd8722971, 24'd8973284, 24'd9107891, 24'd9100153, 24'd8951602, 24'd8691634, 24'd8371699, 24'd8055109, 24'd7804519, 24'd7669518, 
24'd7676824, 24'd7824990, 24'd8084696, 24'd8404545, 24'd8721240, 24'd8972107, 24'd9107501, 24'd9100628, 24'd8952847, 24'd8693404, 24'd8373642, 24'd8056842, 24'd7805698, 24'd7669910, 24'd7676352, 24'd7823747, 24'd8082928, 24'd8402601, 24'd8719506, 24'd8970926, 24'd9107107, 24'd9101097, 24'd8954088, 24'd8695171, 24'd8375585, 24'd8058577, 24'd7806881, 24'd7670308, 24'd7675885, 24'd7822508, 
24'd8081162, 24'd8400658, 24'd8717770, 24'd8969741, 24'd9106707, 24'd9101562, 24'd8955325, 24'd8696936, 24'd8377529, 24'd8060314, 24'd7808068, 24'd7670710, 24'd7675423, 24'd7821273, 24'd8079398, 24'd8398715, 24'd8716031, 24'd8968552, 24'd9106302, 24'd9102022, 24'd8956558, 24'd8698698, 24'd8379472, 24'd8062054, 24'd7809260, 24'd7671118, 24'd7674965, 24'd7820042, 24'd8077636, 24'd8396771, 
24'd8714291, 24'd8967358, 24'd9105892, 24'd9102476, 24'd8957787, 24'd8700459, 24'd8381415, 24'd8063795, 24'd7810455, 24'd7671530, 24'd7674513, 24'd7818815, 24'd8075877, 24'd8394828, 24'd8712548, 24'd8966161, 24'd9105477, 24'd9102926, 24'd8959012, 24'd8702217, 24'd8383359, 24'd8065539, 24'd7811655, 24'd7671948, 24'd7674066, 24'd7817591, 24'd8074120, 24'd8392884, 24'd8710803, 24'd8964959, 
24'd9105057, 24'd9103370, 24'd8960234, 24'd8703973, 24'd8385302, 24'd8067286, 24'd7812858, 24'd7672370, 24'd7673624, 24'd7816372, 24'd8072365, 24'd8390941, 24'd8709055, 24'd8963754, 24'd9104632, 24'd9103810, 24'd8961451, 24'd8705727, 24'd8387246, 24'd8069034, 24'd7814066, 24'd7672798, 24'd7673187, 24'd7815157, 24'd8070612, 24'd8388997, 24'd8707306, 24'd8962544, 24'd9104202, 24'd9104245, 
24'd8962664, 24'd8707479, 24'd8389190, 24'd8070785, 24'd7815277, 24'd7673230, 24'd7672755, 24'd7813946, 24'd8068861, 24'd8387054, 24'd8705554, 24'd8961331, 24'd9103767, 24'd9104674, 24'd8963873, 24'd8709228, 24'd8391133, 24'd8072538, 24'd7816493, 24'd7673668, 24'd7672328, 24'd7812739, 24'd8067113, 24'd8385110, 24'd8703799, 24'd8960113, 24'd9103327, 24'd9105099, 24'd8965078, 24'd8710976, 
24'd8393077, 24'd8074293, 24'd7817712, 24'd7674110, 24'd7671906, 24'd7811536, 24'd8065367, 24'd8383167, 24'd8702043, 24'd8958891, 24'd9102882, 24'd9105518, 24'd8966279, 24'd8712721, 24'd8395020, 24'd8076051, 24'd7818936, 24'd7674558, 24'd7671489, 24'd7810337, 24'd8063623, 24'd8381223, 24'd8700285, 24'd8957666, 24'd9102431, 24'd9105933, 24'd8967476, 24'd8714463, 24'd8396964, 24'd8077811, 
24'd7820164, 24'd7675011, 24'd7671077, 24'd7809142, 24'd8061881, 24'd8379280, 24'd8698524, 24'd8956436, 24'd9101976, 24'd9106342, 24'd8968669, 24'd8716204, 24'd8398907, 24'd8079572, 24'd7821395, 24'd7675468, 24'd7670670, 24'd7807951, 24'd8060142, 24'd8377336, 24'd8696761, 24'd8955203, 24'd9101516, 24'd9106746, 24'd8969858, 24'd8717942, 24'd8400850, 24'd8081336, 24'd7822631, 24'd7675931, 
24'd7670268, 24'd7806764, 24'd8058405, 24'd8375393, 24'd8694996, 24'd8953965, 24'd9101051, 24'd9107146, 24'd8971043, 24'd8719678, 24'd8402794, 24'd8083103, 24'd7823870, 24'd7676398, 24'd7669871, 24'd7805581, 24'd8056670, 24'd8373450, 24'd8693229, 24'd8952724, 24'd9100581, 24'd9107540, 24'd8972224, 24'd8721411, 24'd8404737, 24'd8084871, 24'd7825114, 24'd7676871, 24'd7669480, 24'd7804402, 
24'd8054938, 24'd8371507, 24'd8691459, 24'd8951478, 24'd9100106, 24'd9107930, 24'd8973401, 24'd8723142, 24'd8406680, 24'd8086641, 24'd7826361, 24'd7677348, 24'd7669093, 24'd7803228, 24'd8053208, 24'd8369564, 24'd8689688, 24'd8950229, 24'd9099626, 24'd9108314, 24'd8974573, 24'd8724871, 24'd8408623, 24'd8088414, 24'd7827612, 24'd7677831, 24'd7668711, 24'd7802057, 24'd8051481, 24'd8367621, 
24'd8687914, 24'd8948975, 24'd9099141, 24'd9108693, 24'd8975742, 24'd8726597, 24'd8410566, 24'd8090188, 24'd7828868, 24'd7678319, 24'd7668334, 24'd7800891, 24'd8049755, 24'd8365678, 24'd8686138, 24'd8947718, 24'd9098651, 24'd9109067, 24'd8976906, 24'd8728321, 24'd8412508, 24'd8091965, 24'd7830127, 24'd7678811, 24'd7667963, 24'd7799728, 24'd8048032, 24'd8363735, 24'd8684361, 24'd8946457, 
24'd9098156, 24'd9109436, 24'd8978066, 24'd8730043, 24'd8414451, 24'd8093744, 24'd7831390, 24'd7679309, 24'd7667596, 24'd7798570, 24'd8046312, 24'd8361793, 24'd8682581, 24'd8945192, 24'd9097656, 24'd9109800, 24'd8979222, 24'd8731762, 24'd8416393, 24'd8095525, 24'd7832657, 24'd7679811, 24'd7667235, 24'd7797416, 24'd8044594, 24'd8359851, 24'd8680799, 24'd8943923, 24'd9097151, 24'd9110159, 
24'd8980374, 24'd8733479, 24'd8418335, 24'd8097308, 24'd7833928, 24'd7680319, 24'd7666878, 24'd7796266, 24'd8042878, 24'd8357909, 24'd8679015, 24'd8942650, 24'd9096641, 24'd9110513, 24'd8981522, 24'd8735194, 24'd8420277, 24'd8099093, 24'd7835203, 24'd7680831, 24'd7666527, 24'd7795121, 24'd8041165, 24'd8355967, 24'd8677229, 24'd8941373, 24'd9096126, 24'd9110862, 24'd8982666, 24'd8736906, 
24'd8422219, 24'd8100880, 24'd7836482, 24'd7681348, 24'd7666180, 24'd7793979, 24'd8039454, 24'd8354026, 24'd8675441, 24'd8940092, 24'd9095606, 24'd9111206, 24'd8983805, 24'd8738615, 24'd8424160, 24'd8102669, 24'd7837764, 24'd7681871, 24'd7665839, 24'd7792842, 24'd8037746, 24'd8352084, 24'd8673651, 24'd8938808, 24'd9095081, 24'd9111545, 24'd8984940, 24'd8740323, 24'd8426101, 24'd8104460, 
24'd7839051, 24'd7682398, 24'd7665503, 24'd7791709, 24'd8036040, 24'd8350143, 24'd8671859, 24'd8937519, 24'd9094551, 24'd9111878, 24'd8986071, 24'd8742027, 24'd8428042, 24'd8106253, 24'd7840341, 24'd7682930, 24'd7665172, 24'd7790580, 24'd8034336, 24'd8348202, 24'd8670065, 24'd8936227, 24'd9094017, 24'd9112207, 24'd8987198, 24'd8743730, 24'd8429983, 24'd8108048, 24'd7841635, 24'd7683468, 
24'd7664846, 24'd7789455, 24'd8032635, 24'd8346262, 24'd8668269, 24'd8934931, 24'd9093477, 24'd9112531, 24'd8988321, 24'd8745429, 24'd8431923, 24'd8109845, 24'd7842933, 24'd7684010, 24'd7664525, 24'd7788334, 24'd8030937, 24'd8344322, 24'd8666471, 24'd8933631, 24'd9092932, 24'd9112849, 24'd8989440, 24'd8747126, 24'd8433863, 24'd8111644, 24'd7844235, 24'd7684557, 24'd7664209, 24'd7787218, 
24'd8029241, 24'd8342382, 24'd8664671, 24'd8932328, 24'd9092383, 24'd9113162, 24'd8990554, 24'd8748821, 24'd8435803, 24'd8113445, 24'd7845541, 24'd7685109, 24'd7663898, 24'd7786106, 24'd8027547, 24'd8340442, 24'd8662869, 24'd8931020, 24'd9091828, 24'd9113471, 24'd8991664, 24'd8750513, 24'd8437742, 24'd8115248, 24'd7846850, 24'd7685666, 24'd7663592, 24'd7784998, 24'd8025857, 24'd8338503, 
24'd8661065, 24'd8929709, 24'd9091269, 24'd9113774, 24'd8992770, 24'd8752203, 24'd8439681, 24'd8117052, 24'd7848163, 24'd7686228, 24'd7663291, 24'd7783894, 24'd8024168, 24'd8336564, 24'd8659260, 24'd8928393, 24'd9090705, 24'd9114072, 24'd8993871, 24'd8753890, 24'd8441620, 24'd8118859, 24'd7849481, 24'd7686794, 24'd7662996, 24'd7782794, 24'd8022482, 24'd8334626, 24'd8657452, 24'd8927075, 
24'd9090135, 24'd9114365, 24'd8994969, 24'd8755575, 24'd8443558, 24'd8120667, 24'd7850801, 24'd7687366, 24'd7662705, 24'd7781699, 24'd8020799, 24'd8332688, 24'd8655643, 24'd8925752, 24'd9089561, 24'd9114653, 24'd8996062, 24'd8757257, 24'd8445496, 24'd8122478, 24'd7852126, 24'd7687943, 24'd7662420, 24'd7780608, 24'd8019118, 24'd8330750, 24'd8653831, 24'd8924425, 24'd9088982, 24'd9114936, 
24'd8997151, 24'd8758936, 24'd8447434, 24'd8124290, 24'd7853454, 24'd7688524, 24'd7662140, 24'd7779521, 24'd8017440, 24'd8328813, 24'd8652018, 24'd8923095, 24'd9088398, 24'd9115214, 24'd8998235, 24'd8760613, 24'd8449371, 24'd8126104, 24'd7854786, 24'd7689111, 24'd7661864, 24'd7778439, 24'd8015765, 24'd8326876, 24'd8650203, 24'd8921761, 24'd9087809, 24'd9115486, 24'd8999316, 24'd8762287, 
24'd8451308, 24'd8127920, 24'd7856122, 24'd7689702, 24'd7661594, 24'd7777361, 24'd8014092, 24'd8324939, 24'd8648386, 24'd8920423, 24'd9087215, 24'd9115754, 24'd9000392, 24'd8763958, 24'd8453244, 24'd8129738, 24'd7857462, 24'd7690298, 24'd7661329, 24'd7776287, 24'd8012422, 24'd8323003, 24'd8646568, 24'd8919082, 24'd9086617, 24'd9116016, 24'd9001463, 24'd8765627, 24'd8455180, 24'd8131557, 
24'd7858805, 24'd7690900, 24'd7661069, 24'd7775217, 24'd8010754, 24'd8321068, 24'd8644747, 24'd8917737, 24'd9086013, 24'd9116274, 24'd9002531, 24'd8767294, 24'd8457115, 24'd8133379, 24'd7860152, 24'd7691506, 24'd7660814, 24'd7774152, 24'd8009089, 24'd8319133, 24'd8642925, 24'd8916388, 24'd9085405, 24'd9116526, 24'd9003594, 24'd8768957, 24'd8459050, 24'd8135202, 24'd7861503, 24'd7692117, 
24'd7660565, 24'd7773091, 24'd8007427, 24'd8317198, 24'd8641101, 24'd8915035, 24'd9084791, 24'd9116773, 24'd9004653, 24'd8770618, 24'd8460984, 24'd8137027, 24'd7862857, 24'd7692732, 24'd7660320, 24'd7772034, 24'd8005767, 24'd8315264, 24'd8639275, 24'd8913679, 24'd9084173, 24'd9117015, 24'd9005707, 24'd8772276, 24'd8462918, 24'd8138854, 24'd7864215, 24'd7693353, 24'd7660080, 24'd7770982, 
24'd8004111, 24'd8313330, 24'd8637447, 24'd8912319, 24'd9083550, 24'd9117252, 24'd9006758, 24'd8773932, 24'd8464851, 24'd8140682, 24'd7865577, 24'd7693979, 24'd7659846, 24'd7769934, 24'd8002456, 24'd8311397, 24'd8635618, 24'd8910956, 24'd9082922, 24'd9117484, 24'd9007803, 24'd8775585, 24'd8466784, 24'd8142512, 24'd7866943, 24'd7694609, 24'd7659617, 24'd7768890, 24'd8000805, 24'd8309465, 
24'd8633787, 24'd8909588, 24'd9082289, 24'd9117711, 24'd9008845, 24'd8777235, 24'd8468716, 24'd8144344, 24'd7868312, 24'd7695244, 24'd7659393, 24'd7767851, 24'd7999156, 24'd8307533, 24'd8631954, 24'd8908217, 24'd9081651, 24'd9117933, 24'd9009882, 24'd8778882, 24'd8470648, 24'd8146178, 24'd7869684, 24'd7695885, 24'd7659173, 24'd7766816, 24'd7997510, 24'd8305601, 24'd8630119, 24'd8906843, 
24'd9081008, 24'd9118149, 24'd9010915, 24'd8780527, 24'd8472579, 24'd8148013, 24'd7871061, 24'd7696530, 24'd7658959, 24'd7765785, 24'd7995867, 24'd8303670, 24'd8628283, 24'd8905465, 24'd9080361, 24'd9118361, 24'd9011943, 24'd8782169, 24'd8474510, 24'd8149850, 24'd7872441, 24'd7697180, 24'd7658751, 24'd7764759, 24'd7994226, 24'd8301740, 24'd8626445, 24'd8904083, 24'd9079709, 24'd9118567, 
24'd9012967, 24'd8783808, 24'd8476440, 24'd8151689, 24'd7873824, 24'd7697834, 24'd7658547, 24'd7763737, 24'd7992588, 24'd8299811, 24'd8624606, 24'd8902697, 24'd9079052, 24'd9118768, 24'd9013987, 24'd8785445, 24'd8478369, 24'd8153530, 24'd7875212, 24'd7698494, 24'd7658348, 24'd7762720, 24'd7990953, 24'd8297882, 24'd8622765, 24'd8901308, 24'd9078390, 24'd9118964, 24'd9015002, 24'd8787078, 
24'd8480298, 24'd8155372, 24'd7876602, 24'd7699158, 24'd7658155, 24'd7761707, 24'd7989321, 24'd8295953, 24'd8620922, 24'd8899916, 24'd9077723, 24'd9119155, 24'd9016013, 24'd8788709, 24'd8482226, 24'd8157215, 24'd7877997, 24'd7699828, 24'd7657966, 24'd7760698, 24'd7987691, 24'd8294026, 24'd8619077, 24'd8898520, 24'd9077051, 24'd9119341, 24'd9017020, 24'd8790337, 24'd8484153, 24'd8159061, 
24'd7879395, 24'd7700502, 24'd7657783, 24'd7759694, 24'd7986065, 24'd8292099, 24'd8617231, 24'd8897120, 24'd9076375, 24'd9119522, 24'd9018022, 24'd8791962, 24'd8486080, 24'd8160907, 24'd7880797, 24'd7701181, 24'd7657605, 24'd7758694, 24'd7984441, 24'd8290172, 24'd8615384, 24'd8895716, 24'd9075693, 24'd9119697, 24'd9019020, 24'd8793585, 24'd8488006, 24'd8162756, 24'd7882202, 24'd7701864, 
24'd7657432, 24'd7757698, 24'd7982820, 24'd8288247, 24'd8613534, 24'd8894309, 24'd9075007, 24'd9119868, 24'd9020013, 24'd8795204, 24'd8489931, 24'd8164606, 24'd7883610, 24'd7702553, 24'd7657264, 24'd7756707, 24'd7981202, 24'd8286322, 24'd8611683, 24'd8892899, 24'd9074316, 24'd9120033, 24'd9021002, 24'd8796821, 24'd8491856, 24'd8166458, 24'd7885023, 24'd7703246, 24'd7657101, 24'd7755720, 
24'd7979587, 24'd8284397, 24'd8609831, 24'd8891485, 24'd9073620, 24'd9120193, 24'd9021986, 24'd8798435, 24'd8493780, 24'd8168311, 24'd7886438, 24'd7703944, 24'd7656944, 24'd7754738, 24'd7977974, 24'd8282474, 24'd8607977, 24'd8890067, 24'd9072920, 24'd9120348, 24'd9022966, 24'd8800046, 24'd8495703, 24'd8170166, 24'd7887858, 24'd7704647, 24'd7656791, 24'd7753760, 24'd7976365, 24'd8280551, 
24'd8606122, 24'd8888646, 24'd9072214, 24'd9120498, 24'd9023942, 24'd8801654, 24'd8497625, 24'd8172022, 24'd7889280, 24'd7705355, 24'd7656644, 24'd7752787, 24'd7974758, 24'd8278629, 24'd8604264, 24'd8887222, 24'd9071504, 24'd9120643, 24'd9024913, 24'd8803259, 24'd8499547, 24'd8173880, 24'd7890707, 24'd7706068, 24'd7656502, 24'd7751818, 24'd7973154, 24'd8276708, 24'd8602406, 24'd8885794, 
24'd9070789, 24'd9120782, 24'd9025879, 24'd8804861, 24'd8501468, 24'd8175739, 24'd7892137, 24'd7706785, 24'd7656365, 24'd7750854, 24'd7971553, 24'd8274787, 24'd8600546, 24'd8884362, 24'd9070070, 24'd9120917, 24'd9026842, 24'd8806461, 24'd8503388, 24'd8177600, 24'd7893570, 24'd7707507, 24'd7656233, 24'd7749894, 24'd7969956, 24'd8272868, 24'd8598684, 24'd8882927, 24'd9069345, 24'd9121046, 
24'd9027799, 24'd8808057, 24'd8505307, 24'd8179462, 24'd7895007, 24'd7708234, 24'd7656106, 24'd7748939, 24'd7968361, 24'd8270949, 24'd8596821, 24'd8881489, 24'd9068616, 24'd9121171, 24'd9028752, 24'd8809651, 24'd8507225, 24'd8181326, 24'd7896447, 24'd7708966, 24'd7655984, 24'd7747988, 24'd7966769, 24'd8269031, 24'd8594957, 24'd8880047, 24'd9067882, 24'd9121290, 24'd9029701, 24'd8811241, 
24'd8509143, 24'd8183191, 24'd7897890, 24'd7709702, 24'd7655868, 24'd7747041, 24'd7965180, 24'd8267114, 24'd8593091, 24'd8878601, 24'd9067143, 24'd9121404, 24'd9030645, 24'd8812829, 24'd8511060, 24'd8185058, 24'd7899338, 24'd7710443, 24'd7655756, 24'd7746099, 24'd7963593, 24'd8265197, 24'd8591224, 24'd8877153, 24'd9066400, 24'd9121513, 24'd9031585, 24'd8814413, 24'd8512976, 24'd8186926, 
24'd7900788, 24'd7711189, 24'd7655650, 24'd7745162, 24'd7962010, 24'd8263282, 24'd8589355, 24'd8875700, 24'd9065651, 24'd9121616, 24'd9032520, 24'd8815995, 24'd8514891, 24'd8188795, 24'd7902242, 24'd7711940, 24'd7655549, 24'd7744229, 24'd7960430, 24'd8261367, 24'd8587485, 24'd8874245, 24'd9064898, 24'd9121715, 24'd9033451, 24'd8817574, 24'd8516805, 24'd8190666, 24'd7903699, 24'd7712695, 
24'd7655453, 24'd7743300, 24'd7958853, 24'd8259453, 24'd8585613, 24'd8872786, 24'd9064140, 24'd9121808, 24'd9034377, 24'd8819149, 24'd8518718, 24'd8192538, 24'd7905160, 24'd7713455, 24'd7655362, 24'd7742377, 24'd7957279, 24'd8257541, 24'd8583740, 24'd8871323, 24'd9063378, 24'd9121897, 24'd9035299, 24'd8820722, 24'd8520630, 24'd8194412, 24'd7906624, 24'd7714220, 24'd7655276, 24'd7741457, 
24'd7955708, 24'd8255629, 24'd8581866, 24'd8869857, 24'd9062611, 24'd9121980, 24'd9036216, 24'd8822291, 24'd8522542, 24'd8196287, 24'd7908092, 24'd7714990, 24'd7655196, 24'd7740542, 24'd7954140, 24'd8253718, 24'd8579990, 24'd8868388, 24'd9061839, 24'd9122058, 24'd9037128, 24'd8823858, 24'd8524452, 24'd8198163, 24'd7909563, 24'd7715764, 24'd7655120, 24'd7739632, 24'd7952575, 24'd8251808, 
24'd8578113, 24'd8866916, 24'd9061062, 24'd9122131, 24'd9038036, 24'd8825421, 24'd8526362, 24'd8200041, 24'd7911037, 24'd7716543, 24'd7655050, 24'd7738726, 24'd7951013, 24'd8249899, 24'd8576235, 24'd8865440, 24'd9060280, 24'd9122198, 24'd9038940, 24'd8826982, 24'd8528270, 24'd8201920, 24'd7912515, 24'd7717327, 24'd7654985, 24'd7737825, 24'd7949454, 24'd8247991, 24'd8574355, 24'd8863960, 
24'd9059494, 24'd9122261, 24'd9039839, 24'd8828539, 24'd8530178, 24'd8203800, 24'd7913995, 24'd7718116, 24'd7654925, 24'd7736928, 24'd7947898, 24'd8246084, 24'd8572474, 24'd8862478, 24'd9058703, 24'd9122318, 24'd9040733, 24'd8830093, 24'd8532085, 24'd8205682, 24'd7915480, 24'd7718909, 24'd7654870, 24'd7736036, 24'd7946346, 24'd8244178, 24'd8570592, 24'd8860992, 24'd9057908, 24'd9122371, 
24'd9041623, 24'd8831645, 24'd8533990, 24'd8207565, 24'd7916967, 24'd7719707, 24'd7654820, 24'd7735149, 24'd7944796, 24'd8242272, 24'd8568708, 24'd8859503, 24'd9057108, 24'd9122418, 24'd9042508, 24'd8833193, 24'd8535895, 24'd8209449, 24'd7918458, 24'd7720509, 24'd7654776, 24'd7734266, 24'd7943249, 24'd8240368, 24'd8566824, 24'd8858010, 24'd9056303, 24'd9122460, 24'd9043389, 24'd8834738, 
24'd8537798, 24'd8211334, 24'd7919952, 24'd7721316, 24'd7654736, 24'd7733388, 24'd7941706, 24'd8238465, 24'd8564938, 24'd8856514, 24'd9055493, 24'd9122497, 24'd9044265, 24'd8836279, 24'd8539701, 24'd8213221, 24'd7921450, 24'd7722128, 24'd7654702, 24'd7732514, 24'd7940166, 24'd8236563, 24'd8563050, 24'd8855015, 24'd9054679, 24'd9122528, 24'd9045136, 24'd8837818, 24'd8541602, 24'd8215109, 
24'd7922951, 24'd7722945, 24'd7654673, 24'd7731645, 24'd7938629, 24'd8234663, 24'd8561162, 24'd8853513, 24'd9053860, 24'd9122555, 24'd9046003, 24'd8839354, 24'd8543503, 24'd8216998, 24'd7924455, 24'd7723766, 24'd7654649, 24'd7730780, 24'd7937095, 24'd8232763, 24'd8559272, 24'd8852007, 24'd9053036, 24'd9122576, 24'd9046865, 24'd8840886, 24'd8545402, 24'd8218888, 24'd7925962, 24'd7724592, 
24'd7654630, 24'd7729921, 24'd7935564, 24'd8230864, 24'd8557381, 24'd8850498, 24'd9052208, 24'd9122592, 24'd9047723, 24'd8842415, 24'd8547300, 24'd8220780, 24'd7927472, 24'd7725423, 24'd7654616, 24'd7729065, 24'd7934036, 24'd8228966, 24'd8555489, 24'd8848986, 24'd9051375, 24'd9122604, 24'd9048576, 24'd8843941, 24'd8549197, 24'd8222672, 24'd7928986, 24'd7726258, 24'd7654608, 24'd7728215, 
24'd7932512, 24'd8227070, 24'd8553596, 24'd8847471, 24'd9050538, 24'd9122610, 24'd9049424, 24'd8845464, 24'd8551093, 24'd8224566, 24'd7930503, 24'd7727098, 24'd7654604, 24'd7727369, 24'd7930991, 24'd8225175, 24'd8551701, 24'd8845952, 24'd9049695, 24'd9122610, 24'd9050268, 24'd8846984, 24'd8552988, 24'd8226461, 24'd7932023, 24'd7727943, 24'd7654606, 24'd7726527, 24'd7929473, 24'd8223280, 
24'd8549806, 24'd8844430, 24'd9048848, 24'd9122606, 24'd9051107, 24'd8848500, 24'd8554881, 24'd8228357, 24'd7933547, 24'd7728792, 24'd7654613, 24'd7725691, 24'd7927958, 24'd8221387, 24'd8547909, 24'd8842905, 24'd9047997, 24'd9122597, 24'd9051941, 24'd8850013, 24'd8556774, 24'd8230255, 24'd7935073, 24'd7729645, 24'd7654625, 24'd7724858, 24'd7926447, 24'd8219495, 24'd8546011, 24'd8841377, 
24'd9047141, 24'd9122582, 24'd9052771, 24'd8851523, 24'd8558665, 24'd8232153, 24'd7936603, 24'd7730504, 24'd7654642, 24'd7724031, 24'd7924938, 24'd8217605, 24'd8544112, 24'd8839846, 24'd9046280, 24'd9122562, 24'd9053596, 24'd8853030, 24'd8560555, 24'd8234052, 24'd7938136, 24'd7731367, 24'd7654665, 24'd7723208, 24'd7923433, 24'd8215715, 24'd8542212, 24'd8838311, 24'd9045415, 24'd9122537, 
24'd9054416, 24'd8854533, 24'd8562444, 24'd8235953, 24'd7939672, 24'd7732235, 24'd7654692, 24'd7722390, 24'd7921931, 24'd8213827, 24'd8540311, 24'd8836774, 24'd9044545, 24'd9122507, 24'd9055232, 24'd8856033, 24'd8564332, 24'd8237855, 24'd7941211, 24'd7733107, 24'd7654725, 24'd7721577, 24'd7920433, 24'd8211940, 24'd8538409, 24'd8835233, 24'd9043670, 24'd9122472, 24'd9056043, 24'd8857530, 
24'd8566218, 24'd8239757, 24'd7942754, 24'd7733984, 24'd7654762, 24'd7720768, 24'd7918938, 24'd8210054, 24'd8536506, 24'd8833689, 24'd9042791, 24'd9122432, 24'd9056850, 24'd8859024, 24'd8568103, 24'd8241661, 24'd7944299, 24'd7734865, 24'd7654805, 24'd7719964, 24'd7917446, 24'd8208170, 24'd8534602, 24'd8832142, 24'd9041908, 24'd9122386, 24'd9057651, 24'd8860514, 24'd8569987, 24'd8243566, 
24'd7945848, 24'd7735751, 24'd7654853, 24'd7719164, 24'd7915957, 24'd8206286, 24'd8532696, 24'd8830592, 24'd9041019, 24'd9122336, 24'd9058449, 24'd8862001, 24'd8571870, 24'd8245472, 24'd7947399, 24'd7736642, 24'd7654907, 24'd7718370, 24'd7914472, 24'd8204404, 24'd8530790, 24'd8829039, 24'd9040126, 24'd9122280, 24'd9059241, 24'd8863485, 24'd8573751, 24'd8247378, 24'd7948954, 24'd7737537, 
24'd7654965, 24'd7717580, 24'd7912990, 24'd8202523, 24'd8528883, 24'd8827482, 24'd9039229, 24'd9122219, 24'd9060029, 24'd8864965, 24'd8575631, 24'd8249286, 24'd7950512, 24'd7738436, 24'd7655028, 24'd7716794, 24'd7911511, 24'd8200644, 24'd8526975, 24'd8825923, 24'd9038327, 24'd9122153, 24'd9060811, 24'd8866442, 24'd8577510, 24'd8251195, 24'd7952073, 24'd7739341, 24'd7655097, 24'd7716014, 
24'd7910036, 24'd8198766, 24'd8525066, 24'd8824360, 24'd9037420, 24'd9122082, 24'd9061590, 24'd8867916, 24'd8579388, 24'd8253104, 24'd7953637, 24'd7740250, 24'd7655171, 24'd7715238, 24'd7908564, 24'd8196889, 24'd8523155, 24'd8822795, 24'd9036509, 24'd9122005, 24'd9062363, 24'd8869386, 24'd8581264, 24'd8255015, 24'd7955204, 24'd7741163, 24'd7655250, 24'd7714467, 24'd7907095, 24'd8195014, 
24'd8521244, 24'd8821226, 24'd9035594, 24'd9121924, 24'd9063132, 24'd8870853, 24'd8583139, 24'd8256927, 24'd7956774, 24'd7742081, 24'd7655334, 24'd7713700, 24'd7905630, 24'd8193140, 24'd8519332, 24'd8819655, 24'd9034674, 24'd9121837, 24'd9063896, 24'd8872317, 24'd8585012, 24'd8258839, 24'd7958347, 24'd7743003, 24'd7655423, 24'd7712939, 24'd7904168, 24'd8191267, 24'd8517419, 24'd8818080, 
24'd9033749, 24'd9121745, 24'd9064655, 24'd8873777, 24'd8586884, 24'd8260753, 24'd7959924, 24'd7743930, 24'd7655517, 24'd7712182, 24'd7902710, 24'd8189396, 24'd8515505, 24'd8816502, 24'd9032820, 24'd9121648, 24'd9065410, 24'd8875233, 24'd8588755, 24'd8262667, 24'd7961503, 24'd7744862, 24'd7655617, 24'd7711430, 24'd7901254, 24'd8187526, 24'd8513591, 24'd8814922, 24'd9031886, 24'd9121546, 
24'd9066160, 24'd8876687, 24'd8590624, 24'd8264582, 24'd7963085, 24'd7745798, 24'd7655722, 24'd7710682, 24'd7899803, 24'd8185657, 24'd8511675, 24'd8813338, 24'd9030948, 24'd9121439, 24'd9066905, 24'd8878137, 24'd8592492, 24'd8266498, 24'd7964670, 24'd7746738, 24'd7655831, 24'd7709939, 24'd7898355, 24'd8183790, 24'd8509758, 24'd8811751, 24'd9030005, 24'd9121327, 24'd9067645, 24'd8879583, 
24'd8594358, 24'd8268415, 24'd7966258, 24'd7747683, 24'd7655946, 24'd7709201, 24'd7896910, 24'd8181924, 24'd8507841, 24'd8810162, 24'd9029058, 24'd9121209, 24'd9068381, 24'd8881026, 24'd8596223, 24'd8270333, 24'd7967849, 24'd7748633, 24'd7656066, 24'd7708468, 24'd7895469, 24'd8180060, 24'd8505923, 24'd8808569, 24'd9028106, 24'd9121087, 24'd9069112, 24'd8882466, 24'd8598086, 24'd8272251, 
24'd7969443, 24'd7749587, 24'd7656191, 24'd7707740, 24'd7894031, 24'd8178197, 24'd8504004, 24'd8806974, 24'd9027150, 24'd9120959, 24'd9069838, 24'd8883902, 24'd8599948, 24'd8274171, 24'd7971040, 24'd7750545, 24'd7656322, 24'd7707016, 24'd7892596, 24'd8176336, 24'd8502084, 24'd8805375, 24'd9026189, 24'd9120826, 24'd9070559, 24'd8885335, 24'd8601809, 24'd8276091, 24'd7972640, 24'd7751508, 
24'd7656457, 24'd7706297, 24'd7891165, 24'd8174476, 24'd8500164, 24'd8803774, 24'd9025224, 24'd9120688, 24'd9071275, 24'd8886764, 24'd8603668, 24'd8278012, 24'd7974243, 24'd7752476, 24'd7656598, 24'd7705583, 24'd7889738, 24'd8172618, 24'd8498242, 24'd8802170, 24'd9024254, 24'd9120545, 24'd9071987, 24'd8888189, 24'd8605525, 24'd8279934, 24'd7975849, 24'd7753447, 24'd7656743, 24'd7704874, 
24'd7888314, 24'd8170761, 24'd8496320, 24'd8800563, 24'd9023280, 24'd9120397, 24'd9072694, 24'd8889612, 24'd8607381, 24'd8281856, 24'd7977457, 24'd7754424, 24'd7656894, 24'd7704169, 24'd7886894, 24'd8168906, 24'd8494397, 24'd8798952, 24'd9022301, 24'd9120243, 24'd9073396, 24'd8891030, 24'd8609236, 24'd8283780, 24'd7979069, 24'd7755405, 24'd7657050, 24'd7703470, 24'd7885477, 24'd8167052, 
24'd8492473, 24'd8797340, 24'd9021318, 24'd9120085, 24'd9074093, 24'd8892445, 24'd8611089, 24'd8285704, 24'd7980683, 24'd7756390, 24'd7657211, 24'd7702775, 24'd7884063, 24'd8165200, 24'd8490549, 24'd8795724, 24'd9020331, 24'd9119921, 24'd9074786, 24'd8893857, 24'd8612940, 24'd8287628, 24'd7982300, 24'd7757379, 24'd7657378, 24'd7702085, 24'd7882654, 24'd8163350, 24'd8488624, 24'd8794105, 
24'd9019339, 24'd9119752, 24'd9075473, 24'd8895265, 24'd8614790, 24'd8289554, 24'd7983920, 24'd7758374, 24'd7657549, 24'd7701400, 24'd7881247, 24'd8161501, 24'd8486698, 24'd8792484, 24'd9018343, 24'd9119578, 24'd9076156, 24'd8896670, 24'd8616638, 24'd8291480, 24'd7985543, 24'd7759372, 24'd7657725, 24'd7700719, 24'd7879845, 24'd8159653, 24'd8484772, 24'd8790859, 24'd9017342, 24'd9119399, 
24'd9076834, 24'd8898070, 24'd8618485, 24'd8293407, 24'd7987169, 24'd7760375, 24'd7657907, 24'd7700043, 24'd7878445, 24'd8157807, 24'd8482844, 24'd8789232, 24'd9016337, 24'd9119215, 24'd9077508, 24'd8899468, 24'd8620330, 24'd8295334, 24'd7988797, 24'd7761382, 24'd7658094, 24'd7699373, 24'd7877050, 24'd8155963, 24'd8480917, 24'd8787602, 24'd9015327, 24'd9119026, 24'd9078176, 24'd8900862, 
24'd8622173, 24'd8297262, 24'd7990429, 24'd7762394, 24'd7658286, 24'd7698707, 24'd7875658, 24'd8154121, 24'd8478988, 24'd8785969, 24'd9014314, 24'd9118832, 24'd9078840, 24'd8902252, 24'd8624015, 24'd8299191, 24'd7992063, 24'd7763410, 24'd7658483, 24'd7698046, 24'd7874269, 24'd8152280, 24'd8477059, 24'd8784334, 24'd9013295, 24'd9118632, 24'd9079498, 24'd8903638, 24'd8625855, 24'd8301121, 
24'd7993700, 24'd7764431, 24'd7658685, 24'd7697389, 24'd7872885, 24'd8150441, 24'd8475129, 24'd8782696, 24'd9012273, 24'd9118427, 24'd9080152, 24'd8905021, 24'd8627693, 24'd8303051, 24'd7995340, 24'd7765455, 24'd7658892, 24'd7696738, 24'd7871503, 24'd8148603, 24'd8473199, 24'd8781055, 24'd9011246, 24'd9118218, 24'd9080801, 24'd8906401, 24'd8629530, 24'd8304981, 24'd7996982, 24'd7766485, 
24'd7659104, 24'd7696091, 24'd7870126, 24'd8146767, 24'd8471268, 24'd8779411, 24'd9010214, 24'd9118003, 24'd9081445, 24'd8907777, 24'd8631365, 24'd8306913, 24'd7998627, 24'd7767518, 24'd7659322, 24'd7695449, 24'd7868752, 24'd8144933, 24'd8469337, 24'd8777764, 24'd9009178, 24'd9117783, 24'd9082085, 24'd8909149, 24'd8633199, 24'd8308844, 24'd8000275, 24'd7768556, 24'd7659544, 24'd7694813, 
24'd7867382, 24'd8143100, 24'd8467405, 24'd8776115, 24'd9008138, 24'd9117558, 24'd9082719, 24'd8910517, 24'd8635030, 24'd8310777, 24'd8001926, 24'd7769598, 24'd7659772, 24'd7694181, 24'd7866015, 24'd8141270, 24'd8465472, 24'd8774463, 24'd9007094, 24'd9117327, 24'd9083349, 24'd8911882, 24'd8636860, 24'd8312710, 24'd8003579, 24'd7770645, 24'd7660005, 24'd7693553, 24'd7864652, 24'd8139441, 
24'd8463539, 24'd8772808, 24'd9006045, 24'd9117092, 24'd9083973, 24'd8913243, 24'd8638688, 24'd8314643, 24'd8005235, 24'd7771696, 24'd7660243, 24'd7692931, 24'd7863293, 24'd8137613, 24'd8461605, 24'd8771151, 24'd9004992, 24'd9116852, 24'd9084593, 24'd8914600, 24'd8640515, 24'd8316577, 24'd8006894, 24'd7772751, 24'd7660486, 24'd7692314, 24'd7861937, 24'd8135788, 24'd8459671, 24'd8769491, 
24'd9003934, 24'd9116606, 24'd9085208, 24'd8915954, 24'd8642339, 24'd8318511, 24'd8008555, 24'd7773811, 24'd7660734, 24'd7691701, 24'd7860585, 24'd8133964, 24'd8457736, 24'd8767828, 24'd9002873, 24'd9116355, 24'd9085818, 24'd8917304, 24'd8644162, 24'd8320446, 24'd8010219, 24'd7774875, 24'd7660987, 24'd7691094, 24'd7859237, 24'd8132142, 24'd8455801, 24'd8766163, 24'd9001807, 24'd9116100, 
24'd9086423, 24'd8918651, 24'd8645983, 24'd8322382, 24'd8011886, 24'd7775943, 24'd7661245, 24'd7690491, 24'd7857893, 24'd8130322, 24'd8453865, 24'd8764494, 24'd9000736, 24'd9115839, 24'd9087024, 24'd8919993, 24'd8647803, 24'd8324318, 24'd8013556, 24'd7777016, 24'd7661509, 24'd7689893, 24'd7856552, 24'd8128504, 24'd8451929, 24'd8762824, 24'd8999662, 24'd9115573, 24'd9087619, 24'd8921332, 
24'd8649620, 24'd8326254, 24'd8015228, 24'd7778092, 24'd7661777, 24'd7689300, 24'd7855215, 24'd8126687, 24'd8449993, 24'd8761150, 24'd8998583, 24'd9115302, 24'd9088210, 24'd8922667, 24'd8651436, 24'd8328191, 24'd8016902, 24'd7779173, 24'd7662051, 24'd7688712, 24'd7853882, 24'd8124872, 24'd8448056, 24'd8759475, 24'd8997499, 24'd9115026, 24'd9088795, 24'd8923999, 24'd8653249, 24'd8330128, 
24'd8018579, 24'd7780259, 24'd7662329, 24'd7688129, 24'd7852552, 24'd8123059, 24'd8446118, 24'd8757796, 24'd8996412, 24'd9114744, 24'd9089376, 24'd8925326, 24'd8655061, 24'd8332066, 24'd8020259, 24'd7781348, 24'd7662613, 24'd7687551, 24'd7851226, 24'd8121248, 24'd8444181, 24'd8756115, 24'd8995320, 24'd9114458, 24'd9089952, 24'd8926650, 24'd8656871, 24'd8334004, 24'd8021942, 24'd7782442, 
24'd7662902, 24'd7686977, 24'd7849904, 24'd8119439, 24'd8442242, 24'd8754431, 24'd8994224, 24'd9114167, 24'd9090522, 24'd8927970, 24'd8658680, 24'd8335942, 24'd8023627, 24'd7783540, 24'd7663196, 24'd7686409, 24'd7848586, 24'd8117632, 24'd8440304, 24'd8752745, 24'd8993124, 24'd9113870, 24'd9091088, 24'd8929287, 24'd8660486, 24'd8337881, 24'd8025314, 24'd7784643, 24'd7663495, 24'd7685846, 
24'd7847271, 24'd8115827, 24'd8438365, 24'd8751056, 24'd8992019, 24'd9113569, 24'd9091649, 24'd8930599, 24'd8662290, 24'd8339820, 24'd8027004, 24'd7785749, 24'd7663799, 24'd7685287, 24'd7845961, 24'd8114023, 24'd8436426, 24'd8749365, 24'd8990911, 24'd9113262, 24'd9092205, 24'd8931908, 24'd8664093, 24'd8341759, 24'd8028697, 24'd7786860, 24'd7664108, 24'd7684733, 24'd7844654, 24'd8112222, 
24'd8434486, 24'd8747671, 24'd8989798, 24'd9112950, 24'd9092757, 24'd8933213, 24'd8665893, 24'd8343699, 24'd8030392, 24'd7787975, 24'd7664423, 24'd7684185, 24'd7843351, 24'd8110422, 24'd8432546, 24'd8745974, 24'd8988681, 24'd9112633, 24'd9093303, 24'd8934514, 24'd8667692, 24'd8345639, 24'd8032090, 24'd7789095, 24'd7664742, 24'd7683641, 24'd7842052, 24'd8108625, 24'd8430606, 24'd8744276, 
24'd8987559, 24'd9112311, 24'd9093844, 24'd8935812, 24'd8669488, 24'd8347579, 24'd8033790, 24'd7790218, 24'd7665066, 24'd7683102, 24'd7840756, 24'd8106829, 24'd8428665, 24'd8742574, 24'd8986434, 24'd9111984, 24'd9094380, 24'd8937105, 24'd8671283, 24'd8349520, 24'd8035493, 24'd7791346, 24'd7665396, 24'd7682568, 24'd7839465, 24'd8105035, 24'd8426724, 24'd8740870, 24'd8985304, 24'd9111652, 
24'd9094912, 24'd8938395, 24'd8673076, 24'd8351461, 24'd8037198, 24'd7792478, 24'd7665731, 24'd7682040, 24'd7838177, 24'd8103244, 24'd8424783, 24'd8739164, 24'd8984170, 24'd9111315, 24'd9095438, 24'd8939680, 24'd8674866, 24'd8353402, 24'd8038905, 24'd7793614, 24'd7666070, 24'd7681516, 24'd7836893, 24'd8101454, 24'd8422842, 24'd8737455, 24'd8983032, 24'd9110973, 24'd9095960, 24'd8940962, 
24'd8676655, 24'd8355344, 24'd8040615, 24'd7794754, 24'd7666415, 24'd7680997, 24'd7835613, 24'd8099666, 24'd8420900, 24'd8735744, 24'd8981890, 24'd9110626, 24'd9096476, 24'd8942240, 24'd8678442, 24'd8357285, 24'd8042328, 24'd7795898, 24'd7666765, 24'd7680483, 24'd7834337, 24'd8097881, 24'd8418959, 24'd8734030, 24'd8980743, 24'd9110274, 24'd9096988, 24'd8943514, 24'd8680226, 24'd8359227, 
24'd8044043, 24'd7797047, 24'd7667120, 24'd7679974, 24'd7833065, 24'd8096097, 24'd8417017, 24'd8732314, 24'd8979592, 24'd9109916, 24'd9097494, 24'd8944785, 24'd8682009, 24'd8361170, 24'd8045760, 24'd7798199, 24'd7667479, 24'd7679469, 24'd7831797, 24'd8094316, 24'd8415074, 24'd8730595, 24'd8978438, 24'd9109554, 24'd9097996, 24'd8946051, 24'd8683789, 24'd8363112, 24'd8047480, 24'd7799356, 
24'd7667844, 24'd7678970, 24'd7830532, 24'd8092536, 24'd8413132, 24'd8728875, 24'd8977279, 24'd9109186, 24'd9098492, 24'd8947314, 24'd8685568, 24'd8365054, 24'd8049202, 24'd7800517, 24'd7668214, 24'd7678476, 24'd7829272, 24'd8090759, 24'd8411189, 24'd8727151, 24'd8976116, 24'd9108814, 24'd9098984, 24'd8948572, 24'd8687344, 24'd8366997, 24'd8050926, 24'd7801682, 24'd7668590, 24'd7677987, 
24'd7828015, 24'd8088983, 24'd8409247, 24'd8725426, 24'd8974949, 24'd9108436, 24'd9099471, 24'd8949827, 24'd8689119, 24'd8368940, 24'd8052653, 24'd7802851, 24'd7668970, 24'd7677503, 24'd7826762, 24'd8087210, 24'd8407304, 24'd8723697, 24'd8973777, 24'd9108053, 24'd9099952, 24'd8951077, 24'd8690891, 24'd8370883, 24'd8054382, 24'd7804025, 24'd7669355, 24'd7677024, 24'd7825514, 24'd8085439, 
24'd8405361, 24'd8721967, 24'd8972602, 24'd9107666, 24'd9100429, 24'd8952324, 24'd8692661, 24'd8372826, 24'd8056114, 24'd7805202, 24'd7669745, 24'd7676550, 24'd7824269, 24'd8083670, 24'd8403418, 24'd8720234, 24'd8971423, 24'd9107273, 24'd9100901, 24'd8953567, 24'd8694429, 24'd8374769, 24'd8057848, 24'd7806384, 24'd7670140, 24'd7676080, 24'd7823028, 24'd8081903, 24'd8401474, 24'd8718499, 
24'd8970239, 24'd9106875, 24'd9101367, 24'd8954806, 24'd8696194, 24'd8376712, 24'd8059584, 24'd7807569, 24'd7670541, 24'd7675616, 24'd7821791, 24'd8080138, 24'd8399531, 24'd8716762, 24'd8969052, 24'd9106472, 24'd9101829, 24'd8956041, 24'd8697958, 24'd8378656, 24'd8061323, 24'd7808759, 24'd7670946, 24'd7675157, 24'd7820558, 24'd8078376, 24'd8397588, 24'd8715022, 24'd8967860, 24'd9106065, 
24'd9102286, 24'd8957271, 24'd8699719, 24'd8380599, 24'd8063063, 24'd7809952, 24'd7671356, 24'd7674703, 24'd7819330, 24'd8076616, 24'd8395644, 24'd8713280, 24'd8966664, 24'd9105652, 24'd9102738, 24'd8958498, 24'd8701479, 24'd8382543, 24'd8064807, 24'd7811150, 24'd7671772, 24'd7674253, 24'd7818105, 24'd8074857, 24'd8393701, 24'd8711536, 24'd8965464, 24'd9105234, 24'd9103184, 24'd8959721, 
24'd8703236, 24'd8384486, 24'd8066552, 24'd7812352, 24'd7672192, 24'd7673809, 24'd7816884, 24'd8073101, 24'd8391757, 24'd8709790, 24'd8964261, 24'd9104811, 24'd9103626, 24'd8960940, 24'd8704991, 24'd8386430, 24'd8068300, 24'd7813558, 24'd7672617, 24'd7673370, 24'd7815667, 24'd8071348, 24'd8389814, 24'd8708041, 24'd8963053, 24'd9104383, 24'd9104063, 24'd8962155, 24'd8706743, 24'd8388373, 
24'd8070049, 24'd7814768, 24'd7673048, 24'd7672936, 24'd7814454, 24'd8069596, 24'd8387870, 24'd8706290, 24'd8961841, 24'd9103950, 24'd9104494, 24'd8963366, 24'd8708494, 24'd8390317, 24'd8071802, 24'd7815982, 24'd7673483, 24'd7672507, 24'd7813245, 24'd8067847, 24'd8385926, 24'd8704537, 24'd8960625, 24'd9103512, 24'd9104921, 24'd8964573, 24'd8710242, 24'd8392260, 24'd8073556, 24'd7817200, 
24'd7673924, 24'd7672083, 24'd7812040, 24'd8066100, 24'd8383983, 24'd8702781, 24'd8959405, 24'd9103069, 24'd9105343, 24'd8965775, 24'd8711988, 24'd8394204, 24'd8075312, 24'd7818421, 24'd7674369, 24'd7671664, 24'd7810840, 24'd8064355, 24'd8382039, 24'd8701024, 24'd8958181, 24'd9102621, 24'd9105759, 24'd8966974, 24'd8713731, 24'd8396147, 24'd8077071, 24'd7819647, 24'd7674820, 24'd7671249, 
24'd7809643, 24'd8062613, 24'd8380096, 24'd8699264, 24'd8956953, 24'd9102168, 24'd9106171, 24'd8968169, 24'd8715473, 24'd8398091, 24'd8078832, 24'd7820877, 24'd7675275, 24'd7670840, 24'd7808450, 24'd8060872, 24'd8378152, 24'd8697502, 24'd8955721, 24'd9101710, 24'd9106577, 24'd8969359, 24'd8717212, 24'd8400034, 24'd8080595, 24'd7822111, 24'd7675736, 24'd7670436, 24'd7807262, 24'd8059134, 
24'd8376209, 24'd8695737, 24'd8954485, 24'd9101247, 24'd9106979, 24'd8970546, 24'd8718949, 24'd8401978, 24'd8082360, 24'd7823349, 24'd7676201, 24'd7670037, 24'd7806077, 24'd8057399, 24'd8374266, 24'd8693971, 24'd8953246, 24'd9100779, 24'd9107375, 24'd8971728, 24'd8720683, 24'd8403921, 24'd8084128, 24'd7824591, 24'd7676672, 24'd7669643, 24'd7804897, 24'd8055665, 24'd8372323, 24'd8692203, 
24'd8952002, 24'd9100306, 24'd9107767, 24'd8972907, 24'd8722415, 24'd8405864, 24'd8085897, 24'd7825837, 24'd7677147, 24'd7669255, 24'd7803721, 24'd8053935, 24'd8370380, 24'd8690432, 24'd8950754, 24'd9099828, 24'd9108153, 24'd8974081, 24'd8724145, 24'd8407807, 24'd8087669, 24'd7827086, 24'd7677628, 24'd7668871, 24'd7802548, 24'd8052206, 24'd8368437, 24'd8688659, 24'd8949502, 24'd9099345, 
24'd9108534, 24'd8975251, 24'd8725873, 24'd8409750, 24'd8089443, 24'd7828340, 24'd7678113, 24'd7668492, 24'd7801380, 24'd8050480, 24'd8366494, 24'd8686885, 24'd8948247, 24'd9098857, 24'd9108911, 24'd8976417, 24'd8727598, 24'd8411692, 24'd8091219, 24'd7829598, 24'd7678604, 24'd7668118, 24'd7800216, 24'd8048756, 24'd8364551, 24'd8685108, 24'd8946987, 24'd9098364, 24'd9109282, 24'd8977579, 
24'd8729320, 24'd8413635, 24'd8092997, 24'd7830859, 24'd7679099, 24'd7667749, 24'd7799056, 24'd8047034, 24'd8362609, 24'd8683329, 24'd8945724, 24'd9097866, 24'd9109648, 24'd8978737, 24'd8731041, 24'd8415577, 24'd8094777, 24'd7832125, 24'd7679599, 24'd7667386, 24'd7797901, 24'd8045315, 24'd8360667, 24'd8681548, 24'd8944456, 24'd9097363, 24'd9110009, 24'd8979891, 24'd8732758, 24'd8417519, 
24'd8096559, 24'd7833394, 24'd7680105, 24'd7667027, 24'd7796749, 24'd8043598, 24'd8358725, 24'd8679765, 24'd8943185, 24'd9096856, 24'd9110365, 24'd8981040, 24'd8734474, 24'd8419461, 24'd8098343, 24'd7834667, 24'd7680615, 24'd7666674, 24'd7795602, 24'd8041884, 24'd8356783, 24'd8677979, 24'd8941910, 24'd9096343, 24'd9110716, 24'd8982186, 24'd8736187, 24'd8421403, 24'd8100129, 24'd7835944, 
24'd7681130, 24'd7666325, 24'd7794458, 24'd8040172, 24'd8354841, 24'd8676192, 24'd8940631, 24'd9095825, 24'd9111062, 24'd8983327, 24'd8737898, 24'd8423345, 24'd8101917, 24'd7837225, 24'd7681651, 24'd7665982, 24'd7793319, 24'd8038463, 24'd8352900, 24'd8674403, 24'd8939348, 24'd9095302, 24'd9111403, 24'd8984464, 24'd8739606, 24'd8425286, 24'd8103707, 24'd7838510, 24'd7682176, 24'd7665643, 
24'd7792184, 24'd8036756, 24'd8350959, 24'd8672612, 24'd8938061, 24'd9094775, 24'd9111739, 24'd8985597, 24'd8741312, 24'd8427227, 24'd8105500, 24'd7839799, 24'd7682706, 24'd7665310, 24'd7791053, 24'd8035051, 24'd8349018, 24'd8670819, 24'd8936771, 24'd9094242, 24'd9112070, 24'd8986725, 24'd8743015, 24'd8429168, 24'd8107294, 24'd7841091, 24'd7683241, 24'd7664982, 24'd7789927, 24'd8033349, 
24'd8347077, 24'd8669023, 24'd8935476, 24'd9093704, 24'd9112395, 24'd8987850, 24'd8744716, 24'd8431108, 24'd8109090, 24'd7842388, 24'd7683781, 24'd7664659, 24'd7788804, 24'd8031650, 24'd8345137, 24'd8667226, 24'd8934178, 24'd9093162, 24'd9112716, 24'd8988970, 24'd8746414, 24'd8433048, 24'd8110888, 24'd7843688, 24'd7684326, 24'd7664341, 24'd7787686, 24'd8029953, 24'd8343197, 24'd8665427, 
24'd8932876, 24'd9092614, 24'd9113031, 24'd8990086, 24'd8748110, 24'd8434988, 24'd8112688, 24'd7844992, 24'd7684876, 24'd7664028, 24'd7786572, 24'd8028258, 24'd8341257, 24'd8663626, 24'd8931570, 24'd9092062, 24'd9113342, 24'd8991198, 24'd8749803, 24'd8436928, 24'd8114490, 24'd7846300, 24'd7685431, 24'd7663720, 24'd7785463, 24'd8026566, 24'd8339318, 24'd8661823, 24'd8930260, 24'd9091505, 
24'd9113647, 24'd8992306, 24'd8751494, 24'd8438867, 24'd8116294, 24'd7847611, 24'd7685991, 24'd7663417, 24'd7784357, 24'd8024877, 24'd8337379, 24'd8660018, 24'd8928946, 24'd9090942, 24'd9113947, 24'd8993409, 24'd8753182, 24'd8440806, 24'd8118100, 24'd7848927, 24'd7686556, 24'd7663119, 24'd7783256, 24'd8023190, 24'd8335440, 24'd8658212, 24'd8927629, 24'd9090375, 24'd9114243, 24'd8994508, 
24'd8754867, 24'd8442744, 24'd8119907, 24'd7850246, 24'd7687125, 24'd7662827, 24'd7782159, 24'd8021506, 24'd8333502, 24'd8656403, 24'd8926308, 24'd9089803, 24'd9114533, 24'd8995603, 24'd8756550, 24'd8444682, 24'd8121717, 24'd7851569, 24'd7687700, 24'd7662539, 24'd7781066, 24'd8019824, 24'd8331564, 24'd8654592, 24'd8924983, 24'd9089226, 24'd9114818, 24'd8996694, 24'd8758231, 24'd8446620, 
24'd8123529, 24'd7852896, 24'd7688279, 24'd7662257, 24'd7779977, 24'd8018145, 24'd8329626, 24'd8652780, 24'd8923654, 24'd9088644, 24'd9115098, 24'd8997780, 24'd8759909, 24'd8448557, 24'd8125342, 24'd7854226, 24'd7688864, 24'd7661979, 24'd7778893, 24'd8016468, 24'd8327689, 24'd8650966, 24'd8922322, 24'd9088057, 24'd9115372, 24'd8998862, 24'd8761584, 24'd8450494, 24'd8127157, 24'd7855561, 
24'd7689453, 24'd7661707, 24'd7777813, 24'd8014794, 24'd8325753, 24'd8649150, 24'd8920986, 24'd9087465, 24'd9115642, 24'd8999940, 24'd8763257, 24'd8452431, 24'd8128974, 24'd7856899, 24'd7690047, 24'd7661440, 24'd7776737, 24'd8013123, 24'd8323816, 24'd8647332, 24'd8919646, 24'd9086869, 24'd9115907, 24'd9001014, 24'd8764927, 24'd8454367, 24'd8130793, 24'd7858240, 24'd7690646, 24'd7661178, 
24'd7775666, 24'd8011454, 24'd8321881, 24'd8645512, 24'd8918302, 24'd9086267, 24'd9116166, 24'd9002083, 24'd8766594, 24'd8456302, 24'd8132614, 24'd7859586, 24'd7691250, 24'd7660921, 24'd7774599, 24'd8009788, 24'd8319945, 24'd8643690, 24'd8916955, 24'd9085661, 24'd9116421, 24'd9003148, 24'd8768259, 24'd8458237, 24'd8134436, 24'd7860935, 24'd7691859, 24'd7660669, 24'd7773536, 24'd8008125, 
24'd8318011, 24'd8641867, 24'd8915604, 24'd9085049, 24'd9116670, 24'd9004209, 24'd8769921, 24'd8460172, 24'd8136260, 24'd7862288, 24'd7692473, 24'd7660422, 24'd7772478, 24'd8006464, 24'd8316076, 24'd8640042, 24'd8914249, 24'd9084433, 24'd9116914, 24'd9005265, 24'd8771580, 24'd8462106, 24'd8138086, 24'd7863644, 24'd7693092, 24'd7660180, 24'd7771424, 24'd8004806, 24'd8314142, 24'd8638215, 
24'd8912891, 24'd9083812, 24'd9117153, 24'd9006317, 24'd8773237, 24'd8464039, 24'd8139914, 24'd7865005, 24'd7693715, 24'd7659944, 24'd7770374, 24'd8003151, 24'd8312209, 24'd8636387, 24'd8911529, 24'd9083186, 24'd9117387, 24'd9007365, 24'd8774891, 24'd8465972, 24'd8141743, 24'd7866369, 24'd7694344, 24'd7659712, 24'd7769328, 24'd8001498, 24'd8310276, 24'd8634556, 24'd8910163, 24'd9082555, 
24'd9117616, 24'd9008408, 24'd8776542, 24'd8467905, 24'd8143575, 24'd7867736, 24'd7694977, 24'd7659486, 24'd7768287, 24'd7999848, 24'd8308344, 24'd8632724, 24'd8908794, 24'd9081920, 24'd9117840, 24'd9009447, 24'd8778191, 24'd8469837, 24'd8145408, 24'd7869107, 24'd7695615, 24'd7659265, 24'd7767250, 24'd7998201, 24'd8306413, 24'd8630890, 24'd8907421, 24'd9081279, 24'd9118059, 24'd9010482, 
24'd8779837, 24'd8471768, 24'd8147242, 24'd7870482, 24'd7696258, 24'd7659049, 24'd7766218, 24'd7996557, 24'd8304481, 24'd8629055, 24'd8906044, 24'd9080634, 24'd9118272, 24'd9011512, 24'd8781480, 24'd8473699, 24'd8149079, 24'd7871861, 24'd7696906, 24'd7658838, 24'd7765190, 24'd7994915, 24'd8302551, 24'd8627218, 24'd8904664, 24'd9079983, 24'd9118481, 24'd9012538, 24'd8783120, 24'd8475629, 
24'd8150917, 24'd7873243, 24'd7697559, 24'd7658632, 24'd7764166, 24'd7993276, 24'd8300621, 24'd8625379, 24'd8903280, 24'd9079328, 24'd9118684, 24'd9013559, 24'd8784758, 24'd8477559, 24'd8152756, 24'd7874628, 24'd7698216, 24'd7658431, 24'd7763147, 24'd7991640, 24'd8298692, 24'd8623538, 24'd8901892, 24'd9078668, 24'd9118882, 24'd9014576, 24'd8786392, 24'd8479488, 24'd8154598, 24'd7876018, 
24'd7698879, 24'd7658235, 24'd7762132, 24'd7990006, 24'd8296763, 24'd8621696, 24'd8900501, 24'd9078003, 24'd9119075, 24'd9015589, 24'd8788024, 24'd8481416, 24'd8156441, 24'd7877411, 24'd7699546, 24'd7658045, 24'd7761121, 24'd7988376, 24'd8294835, 24'd8619852, 24'd8899106, 24'd9077334, 24'd9119263, 24'd9016598, 24'd8789654, 24'd8483343, 24'd8158285, 24'd7878807, 24'd7700218, 24'd7657860, 
24'd7760115, 24'd7986748, 24'd8292908, 24'd8618007, 24'd8897708, 24'd9076659, 24'd9119446, 24'd9017602, 24'd8791280, 24'd8485270, 24'd8160131, 24'd7880207, 24'd7700895, 24'd7657679, 24'd7759113, 24'd7985123, 24'd8290981, 24'd8616160, 24'd8896306, 24'd9075980, 24'd9119624, 24'd9018601, 24'd8792904, 24'd8487197, 24'd8161979, 24'd7881611, 24'd7701576, 24'd7657504, 24'd7758116, 24'd7983501, 
24'd8289055, 24'd8614311, 24'd8894901, 24'd9075296, 24'd9119797, 24'd9019596, 24'd8794524, 24'd8489122, 24'd8163829, 24'd7883018, 24'd7702263, 24'd7657334, 24'd7757123, 24'd7981881, 24'd8287130, 24'd8612461, 24'd8893492, 24'd9074607, 24'd9119964, 24'd9020587, 24'd8796142, 24'd8491047, 24'd8165680, 24'd7884429, 24'd7702954, 24'd7657169, 24'd7756134, 24'd7980265, 24'd8285205, 24'd8610609, 
24'd8892079, 24'd9073913, 24'd9120126, 24'd9021573, 24'd8797757, 24'd8492972, 24'd8167532, 24'd7885843, 24'd7703650, 24'd7657009, 24'd7755150, 24'd7978651, 24'd8283282, 24'd8608756, 24'd8890663, 24'd9073215, 24'd9120284, 24'd9022555, 24'd8799370, 24'd8494895, 24'd8169386, 24'd7887261, 24'd7704351, 24'd7656855, 24'd7754171, 24'd7977040, 24'd8281359, 24'd8606901, 24'd8889244, 24'd9072511, 
24'd9120436, 24'd9023533, 24'd8800979, 24'd8496818, 24'd8171242, 24'd7888682, 24'd7705057, 24'd7656705, 24'd7753195, 24'd7975433, 24'd8279436, 24'd8605045, 24'd8887821, 24'd9071803, 24'd9120583, 24'd9024505, 24'd8802585, 24'd8498740, 24'd8173099, 24'd7890107, 24'd7705768, 24'd7656561, 24'd7752225, 24'd7973828, 24'd8277515, 24'd8603187, 24'd8886394, 24'd9071090, 24'd9120724, 24'd9025474, 
24'd8804189, 24'd8500661, 24'd8174958, 24'd7891536, 24'd7706483, 24'd7656422, 24'd7751258, 24'd7972226, 24'd8275594, 24'd8601327, 24'd8884964, 24'd9070373, 24'd9120861, 24'd9026438, 24'd8805789, 24'd8502581, 24'd8176818, 24'd7892967, 24'd7707203, 24'd7656287, 24'd7750297, 24'd7970626, 24'd8273674, 24'd8599466, 24'd8883530, 24'd9069650, 24'd9120993, 24'd9027398, 24'd8807387, 24'd8504501, 
24'd8178680, 24'd7894403, 24'd7707928, 24'd7656158, 24'd7749339, 24'd7969030, 24'd8271755, 24'd8597604, 24'd8882093, 24'd9068923, 24'd9121119, 24'd9028353, 24'd8808982, 24'd8506420, 24'd8180543, 24'd7895841, 24'd7708658, 24'd7656035, 24'd7748387, 24'd7967437, 24'd8269836, 24'd8595740, 24'd8880653, 24'd9068191, 24'd9121240, 24'd9029303, 24'd8810574, 24'd8508338, 24'd8182407, 24'd7897284, 
24'd7709392, 24'd7655916, 24'd7747438, 24'd7965847, 24'd8267919, 24'd8593875, 24'd8879209, 24'd9067454, 24'd9121356, 24'd9030249, 24'd8812162, 24'd8510255, 24'd8184273, 24'd7898729, 24'd7710131, 24'd7655802, 24'd7746494, 24'd7964259, 24'd8266002, 24'd8592008, 24'd8877762, 24'd9066712, 24'd9121467, 24'd9031191, 24'd8813748, 24'd8512171, 24'd8186141, 24'd7900178, 24'd7710875, 24'd7655694, 
24'd7745555, 24'd7962675, 24'd8264086, 24'd8590140, 24'd8876311, 24'd9065966, 24'd9121573, 24'd9032128, 24'd8815331, 24'd8514086, 24'd8188010, 24'd7901631, 24'd7711624, 24'd7655591, 24'd7744620, 24'd7961094, 24'd8262171, 24'd8588270, 24'd8874857, 24'd9065215, 24'd9121674, 24'd9033061, 24'd8816911, 24'd8516001, 24'd8189880, 24'd7903087, 24'd7712377, 24'd7655492, 24'd7743690, 24'd7959515, 
24'd8260257, 24'd8586399, 24'd8873399, 24'd9064459, 24'd9121770, 24'd9033989, 24'd8818488, 24'd8517915, 24'd8191752, 24'd7904546, 24'd7713135, 24'd7655399, 24'd7742764, 24'd7957940, 24'd8258344, 24'd8584527, 24'd8871938, 24'd9063699, 24'd9121860, 24'd9034912, 24'd8820062, 24'd8519827, 24'd8193625, 24'd7906009, 24'd7713898, 24'd7655312, 24'd7741843, 24'd7956367, 24'd8256432, 24'd8582653, 
24'd8870474, 24'd9062933, 24'd9121945, 24'd9035831, 24'd8821633, 24'd8521739, 24'd8195499, 24'd7907475, 24'd7714666, 24'd7655229, 24'd7740926, 24'd7954798, 24'd8254520, 24'd8580778, 24'd8869006, 24'd9062163, 24'd9122026, 24'd9036746, 24'd8823200, 24'd8523650, 24'd8197375, 24'd7908944, 24'd7715438, 24'd7655151, 24'd7740014, 24'd7953232, 24'd8252610, 24'd8578902, 24'd8867535, 24'd9061389, 
24'd9122101, 24'd9037656, 24'd8824765, 24'd8525560, 24'd8199252, 24'd7910417, 24'd7716215, 24'd7655079, 24'd7739106, 24'd7951669, 24'd8250701, 24'd8577024, 24'd8866060, 24'd9060609, 24'd9122170, 24'd9038561, 24'd8826327, 24'd8527469, 24'd8201130, 24'd7911893, 24'd7716997, 24'd7655012, 24'd7738203, 24'd7950108, 24'd8248792, 24'd8575145, 24'd8864582, 24'd9059825, 24'd9122235, 24'd9039462, 
24'd8827885, 24'd8529377, 24'd8203010, 24'd7913373, 24'd7717784, 24'd7654949, 24'd7737305, 24'd7948551, 24'd8246885, 24'd8573264, 24'd8863101, 24'd9059036, 24'd9122295, 24'd9040358, 24'd8829441, 24'd8531284, 24'd8204891, 24'd7914856, 24'd7718575, 24'd7654892, 24'd7736411, 24'd7946997, 24'd8244978, 24'd8571383, 24'd8861616, 24'd9058243, 24'd9122349, 24'd9041250, 24'd8830993, 24'd8533190, 
24'd8206774, 24'd7916342, 24'd7719371, 24'd7654840, 24'd7735521, 24'd7945446, 24'd8243073, 24'd8569500, 24'd8860129, 24'd9057444, 24'd9122399, 24'd9042137, 24'd8832543, 24'd8535095, 24'd8208657, 24'd7917832, 24'd7720172, 24'd7654794, 24'd7734636, 24'd7943899, 24'd8241168, 24'd8567615, 24'd8858637, 24'd9056641, 24'd9122443, 24'd9043019, 24'd8834089, 24'd8536999, 24'd8210542, 24'd7919324, 
24'd7720977, 24'd7654752, 24'd7733756, 24'd7942354, 24'd8239265, 24'd8565730, 24'd8857143, 24'd9055834, 24'd9122482, 24'd9043897, 24'd8835632, 24'd8538902, 24'd8212428, 24'd7920820, 24'd7721787, 24'd7654716, 24'd7732881, 24'd7940812, 24'd8237362, 24'd8563843, 24'd8855645, 24'd9055021, 24'd9122516, 24'd9044771, 24'd8837172, 24'd8540804, 24'd8214316, 24'd7922320, 24'd7722601, 24'd7654684, 
24'd7732009, 24'd7939274, 24'd8235461, 24'd8561955, 24'd8854144, 24'd9054204, 24'd9122544, 24'd9045639, 24'd8838709, 24'd8542704, 24'd8216204, 24'd7923822, 24'd7723421, 24'd7654658, 24'd7731143, 24'd7937739, 24'd8233561, 24'd8560066, 24'd8852640, 24'd9053383, 24'd9122568, 24'd9046503, 24'd8840243, 24'd8544604, 24'd8218094, 24'd7925328, 24'd7724245, 24'd7654637, 24'd7730281, 24'd7936207, 
24'd8231661, 24'd8558176, 24'd8851132, 24'd9052557, 24'd9122586, 24'd9047363, 24'd8841773, 24'd8546503, 24'd8219985, 24'd7926838, 24'd7725073, 24'd7654621, 24'd7729424, 24'd7934678, 24'd8229763, 24'd8556284, 24'd8849622, 24'd9051726, 24'd9122600, 24'd9048218, 24'd8843301, 24'd8548400, 24'd8221877, 24'd7928350, 24'd7725907, 24'd7654611, 24'd7728571, 24'd7933152, 24'd8227866, 24'd8554391, 
24'd8848108, 24'd9050890, 24'd9122608, 24'd9049068, 24'd8844825, 24'd8550297, 24'd8223771, 24'd7929866, 24'd7726745, 24'd7654605, 24'd7727723, 24'd7931629, 24'd8225971, 24'd8552497, 24'd8846590, 24'd9050050, 24'd9122611, 24'd9049914, 24'd8846346, 24'd8552192, 24'd8225665, 24'd7931384, 24'd7727587, 24'd7654605, 24'd7726880, 24'd7930110, 24'd8224076, 24'd8550602, 24'd8845070, 24'd9049205, 
24'd9122609, 24'd9050755, 24'd8847863, 24'd8554086, 24'd8227561, 24'd7932906, 24'd7728434, 24'd7654609, 24'd7726041, 24'd7928594, 24'd8222182, 24'd8548706, 24'd8843546, 24'd9048355, 24'd9122601, 24'd9051591, 24'd8849378, 24'd8555979, 24'd8229458, 24'd7934432, 24'd7729286, 24'd7654619, 24'd7725207, 24'd7927081, 24'd8220290, 24'd8546809, 24'd8842020, 24'd9047501, 24'd9122589, 24'd9052423, 
24'd8850889, 24'd8557871, 24'd8231355, 24'd7935960, 24'd7730143, 24'd7654634, 24'd7724378, 24'd7925571, 24'd8218399, 24'd8544910, 24'd8840490, 24'd9046642, 24'd9122571, 24'd9053250, 24'd8852397, 24'd8559761, 24'd8233254, 24'd7937492, 24'd7731004, 24'd7654655, 24'd7723553, 24'd7924065, 24'd8216509, 24'd8543011, 24'd8838956, 24'd9045779, 24'd9122548, 24'd9054072, 24'd8853902, 24'd8561651, 
24'd8235155, 24'd7939026, 24'd7731870, 24'd7654680, 24'd7722733, 24'd7922562, 24'd8214620, 24'd8541110, 24'd8837420, 24'd9044911, 24'd9122521, 24'd9054890, 24'd8855404, 24'd8563539, 24'd8237056, 24'd7940564, 24'd7732740, 24'd7654710, 24'd7721918, 24'd7921062, 24'd8212732, 24'd8539208, 24'd8835881, 24'd9044038, 24'd9122488, 24'd9055703, 24'd8856902, 24'd8565426, 24'd8238958, 24'd7942105, 
24'd7733615, 24'd7654746, 24'd7721107, 24'd7919565, 24'd8210846, 24'd8537306, 24'd8834338, 24'd9043161, 24'd9122449, 24'd9056512, 24'd8858397, 24'd8567312, 24'd8240861, 24'd7943650, 24'd7734494, 24'd7654787, 24'd7720301, 24'd7918072, 24'd8208961, 24'd8535402, 24'd8832792, 24'd9042279, 24'd9122406, 24'd9057315, 24'd8859889, 24'd8569196, 24'd8242766, 24'd7945197, 24'd7735378, 24'd7654833, 
24'd7719500, 24'd7916582, 24'd8207077, 24'd8533497, 24'd8831243, 24'd9041393, 24'd9122358, 24'd9058114, 24'd8861377, 24'd8571079, 24'd8244671, 24'd7946747, 24'd7736267, 24'd7654884, 24'd7718703, 24'd7915095, 24'd8205195, 24'd8531591, 24'd8829691, 24'd9040502, 24'd9122304, 24'd9058909, 24'd8862862, 24'd8572961, 24'd8246577, 24'd7948301, 24'd7737160, 24'd7654940, 24'd7717911, 24'd7913612, 
24'd8203313, 24'd8529684, 24'd8828136, 24'd9039606, 24'd9122245, 24'd9059698, 24'd8864344, 24'd8574842, 24'd8248485, 24'd7949857, 24'd7738058, 24'd7655001, 24'd7717124, 24'd7912132, 24'd8201433, 24'd8527776, 24'd8826578, 24'd9038706, 24'd9122181, 24'd9060483, 24'd8865822, 24'd8576721, 24'd8250393, 24'd7951417, 24'd7738960, 24'd7655068, 24'd7716341, 24'd7910655, 24'd8199555, 24'd8525868, 
24'd8825017, 24'd9037802, 24'd9122112, 24'd9061263, 24'd8867297, 24'd8578599, 24'd8252302, 24'd7952980, 24'd7739867, 24'd7655139, 24'd7715563, 24'd7909182, 24'd8197677, 24'd8523958, 24'd8823453, 24'd9036893, 24'd9122038, 24'd9062039, 24'd8868769, 24'd8580476, 24'd8254212, 24'd7954546, 24'd7740779, 24'd7655216, 24'd7714790, 24'd7907712, 24'd8195801, 24'd8522047, 24'd8821885, 24'd9035979, 
24'd9121959, 24'd9062810, 24'd8870237, 24'd8582351, 24'd8256124, 24'd7956114, 24'd7741695, 24'd7655298, 24'd7714022, 24'd7906245, 24'd8193927, 24'd8520135, 24'd8820315, 24'd9035061, 24'd9121874, 24'd9063576, 24'd8871702, 24'd8584225, 24'd8258036, 24'd7957686, 24'd7742615, 24'd7655385, 24'd7713258, 24'd7904782, 24'd8192053, 24'd8518223, 24'd8818742, 24'd9034138, 24'd9121785, 24'd9064337, 
24'd8873164, 24'd8586098, 24'd8259949, 24'd7959261, 24'd7743540, 24'd7655477, 24'd7712499, 24'd7903322, 24'd8190181, 24'd8516309, 24'd8817165, 24'd9033210, 24'd9121690, 24'd9065094, 24'd8874622, 24'd8587969, 24'd8261863, 24'd7960839, 24'd7744470, 24'd7655574, 24'd7711745, 24'd7901865, 24'd8188311, 24'd8514395, 24'd8815586, 24'd9032279, 24'd9121590, 24'd9065845, 24'd8876077, 24'd8589839, 
24'd8263778, 24'd7962420, 24'd7745404, 24'd7655677, 24'd7710995, 24'd7900412, 24'd8186442, 24'd8512480, 24'd8814004, 24'd9031342, 24'd9121485, 24'd9066592, 24'd8877528, 24'd8591707, 24'd8265693, 24'd7964004, 24'd7746343, 24'd7655785, 24'd7710251, 24'd7898963, 24'd8184574, 24'd8510564, 24'd8812418, 24'd9030401, 24'd9121375, 24'd9067335, 24'd8878976, 24'd8593574, 24'd8267610, 24'd7965591, 
24'd7747286, 24'd7655897, 24'd7709511, 24'd7897516, 24'd8182708, 24'd8508647, 24'd8810830, 24'd9029456, 24'd9121259, 24'd9068072, 24'd8880420, 24'd8595440, 24'd8269527, 24'd7967180, 24'd7748233, 24'd7656015, 24'd7708776, 24'd7896074, 24'd8180843, 24'd8506729, 24'd8809238, 24'd9028506, 24'd9121139, 24'd9068805, 24'd8881862, 24'd8597304, 24'd8271445, 24'd7968773, 24'd7749186, 24'd7656138, 
24'd7708045, 24'd7894634, 24'd8178980, 24'd8504810, 24'd8807644, 24'd9027552, 24'd9121013, 24'd9069533, 24'd8883299, 24'd8599166, 24'd8273365, 24'd7970369, 24'd7750142, 24'd7656266, 24'd7707320, 24'd7893198, 24'd8177118, 24'd8502891, 24'd8806047, 24'd9026593, 24'd9120883, 24'd9070256, 24'd8884733, 24'd8601028, 24'd8275284, 24'd7971968, 24'd7751103, 24'd7656400, 24'd7706599, 24'd7891766, 
24'd8175257, 24'd8500970, 24'd8804447, 24'd9025630, 24'd9120747, 24'd9070975, 24'd8886164, 24'd8602887, 24'd8277205, 24'd7973569, 24'd7752069, 24'd7656538, 24'd7705883, 24'd7890337, 24'd8173399, 24'd8499049, 24'd8802844, 24'd9024662, 24'd9120606, 24'd9071689, 24'd8887591, 24'd8604745, 24'd8279127, 24'd7975174, 24'd7753039, 24'd7656682, 24'd7705171, 24'd7888912, 24'd8171541, 24'd8497127, 
24'd8801238, 24'd9023690, 24'd9120460, 24'd9072398, 24'd8889015, 24'd8606602, 24'd8281049, 24'd7976781, 24'd7754013, 24'd7656830, 24'd7704465, 24'd7887490, 24'd8169685, 24'd8495205, 24'd8799629, 24'd9022713, 24'd9120308, 24'd9073102, 24'd8890435, 24'd8608457, 24'd8282972, 24'd7978391, 24'd7754992, 24'd7656984, 24'd7703763, 24'd7886071, 24'd8167831, 24'd8493282, 24'd8798017, 24'd9021732, 
24'd9120152, 24'd9073801, 24'd8891851, 24'd8610311, 24'd8284895, 24'd7980005, 24'd7755975, 24'd7657143, 24'd7703066, 24'd7884657, 24'd8165978, 24'd8491357, 24'd8796403, 24'd9020746, 24'd9119991, 24'd9074495, 24'd8893264, 24'd8612163, 24'd8286820, 24'd7981621, 24'd7756963, 24'd7657307, 24'd7702374, 24'd7883245, 24'd8164127, 24'd8489433, 24'd8794785, 24'd9019756, 24'd9119824, 24'd9075185, 
24'd8894674, 24'd8614013, 24'd8288745, 24'd7983239, 24'd7757955, 24'd7657476, 24'd7701687, 24'd7881838, 24'd8162277, 24'd8487507, 24'd8793165, 24'd9018762, 24'd9119652, 24'd9075870, 24'd8896080, 24'd8615862, 24'd8290671, 24'd7984861, 24'd7758952, 24'd7657651, 24'd7701004, 24'd7880433, 24'd8160429, 24'd8485581, 24'd8791542, 24'd9017763, 24'd9119475, 24'd9076550, 24'd8897482, 24'd8617709, 
24'd8292597, 24'd7986486, 24'd7759953, 24'd7657830, 24'd7700327, 24'd7879033, 24'd8158583, 24'd8483654, 24'd8789916, 24'd9016760, 24'd9119293, 24'd9077225, 24'd8898881, 24'd8619555, 24'd8294525, 24'd7988113, 24'd7760959, 24'd7658015, 24'd7699654, 24'd7877636, 24'd8156738, 24'd8481727, 24'd8788287, 24'd9015752, 24'd9119106, 24'd9077896, 24'd8900277, 24'd8621399, 24'd8296452, 24'd7989743, 
24'd7761968, 24'd7658204, 24'd7698986, 24'd7876242, 24'd8154895, 24'd8479798, 24'd8786656, 24'd9014740, 24'd9118914, 24'd9078561, 24'd8901668, 24'd8623241, 24'd8298381, 24'd7991376, 24'd7762983, 24'd7658399, 24'd7698323, 24'd7874852, 24'd8153053, 24'd8477869, 24'd8785021, 24'd9013724, 24'd9118716, 24'd9079222, 24'd8903056, 24'd8625082, 24'd8300310, 24'd7993012, 24'd7764001, 24'd7658599, 
24'd7697664, 24'd7873466, 24'd8151213, 24'd8475940, 24'd8783384, 24'd9012703, 24'd9118514, 24'd9079878, 24'd8904441, 24'd8626921, 24'd8302240, 24'd7994650, 24'd7765024, 24'd7658804, 24'd7697011, 24'd7872083, 24'd8149375, 24'd8474010, 24'd8781744, 24'd9011677, 24'd9118306, 24'd9080529, 24'd8905822, 24'd8628759, 24'd8304170, 24'd7996292, 24'd7766052, 24'd7659014, 24'd7696362, 24'd7870704, 
24'd8147538, 24'd8472079, 24'd8780102, 24'd9010648, 24'd9118094, 24'd9081175, 24'd8907199, 24'd8630595, 24'd8306101, 24'd7997936, 24'd7767084, 24'd7659230, 24'd7695718, 24'd7869329, 24'd8145703, 24'd8470148, 24'd8778456, 24'd9009614, 24'd9117876, 24'd9081817, 24'd8908573, 24'd8632429, 24'd8308033, 24'd7999583, 24'd7768120, 24'd7659450, 24'd7695079, 24'd7867957, 24'd8143870, 24'd8468216, 
24'd8776808, 24'd9008576, 24'd9117653, 24'd9082453, 24'd8909943, 24'd8634261, 24'd8309965, 24'd8001232, 24'd7769160, 24'd7659676, 24'd7694445, 24'd7866589, 24'd8142038, 24'd8466284, 24'd8775157, 24'd9007533, 24'd9117425, 24'd9083085, 24'd8911309, 24'd8636092, 24'd8311898, 24'd8002884, 24'd7770205, 24'd7659906, 24'd7693816, 24'd7865224, 24'd8140209, 24'd8464351, 24'd8773504, 24'd9006486, 
24'd9117192, 24'd9083712, 24'd8912672, 24'd8637921, 24'd8313831, 24'd8004539, 24'd7771254, 24'd7660142, 24'd7693192, 24'd7863863, 24'd8138381, 24'd8462417, 24'd8771847, 24'd9005435, 24'd9116953, 24'd9084333, 24'd8914031, 24'd8639748, 24'd8315765, 24'd8006197, 24'd7772308, 24'd7660383, 24'd7692572, 24'd7862506, 24'd8136554, 24'd8460483, 24'd8770188, 24'd9004379, 24'd9116710, 24'd9084950, 
24'd8915386, 24'd8641573, 24'd8317699, 24'd8007857, 24'd7773365, 24'd7660629, 24'd7691958, 24'd7861153, 24'd8134730, 24'd8458549, 24'd8768527, 24'd9003319, 24'd9116461, 24'd9085563, 24'd8916738, 24'd8643397, 24'd8319633, 24'd8009520, 24'd7774427, 24'd7660880, 24'd7691348, 24'd7859803, 24'd8132907, 24'd8456614, 24'd8766862, 24'd9002255, 24'd9116208, 24'd9086170, 24'd8918086, 24'd8645219, 
24'd8321569, 24'd8011186, 24'd7775494, 24'd7661136, 24'd7690743, 24'd7858457, 24'd8131086, 24'd8454679, 24'd8765195, 24'd9001186, 24'd9115949, 24'd9086772, 24'd8919430, 24'd8647039, 24'd8323504, 24'd8012854, 24'd7776565, 24'd7661397, 24'd7690144, 24'd7857115, 24'd8129267, 24'd8452743, 24'd8763526, 24'd9000113, 24'd9115685, 24'd9087370, 24'd8920770, 24'd8648857, 24'd8325441, 24'd8014525, 
24'd7777640, 24'd7661664, 24'd7689549, 24'd7855776, 24'd8127450, 24'd8450806, 24'd8761854, 24'd8999036, 24'd9115416, 24'd9087962, 24'd8922107, 24'd8650673, 24'd8327377, 24'd8016198, 24'd7778719, 24'd7661935, 24'd7688958, 24'd7854441, 24'd8125634, 24'd8448869, 24'd8760179, 24'd8997955, 24'd9115142, 24'd9088550, 24'd8923440, 24'd8652488, 24'd8329314, 24'd8017875, 24'd7779802, 24'd7662212, 
24'd7688373, 24'd7853110, 24'd8123821, 24'd8446932, 24'd8758501, 24'd8996869, 24'd9114863, 24'd9089132, 24'd8924769, 24'd8654300, 24'd8331252, 24'd8019553, 24'd7780890, 24'd7662493, 24'd7687793, 24'd7851783, 24'd8122009, 24'd8444995, 24'd8756821, 24'd8995779, 24'd9114579, 24'd9089710, 24'd8926095, 24'd8656111, 24'd8333189, 24'd8021235, 24'd7781982, 24'd7662780, 24'd7687218, 24'd7850459, 
24'd8120199, 24'd8443057, 24'd8755139, 24'd8994685, 24'd9114290, 24'd9090283, 24'd8927416, 24'd8657920, 24'd8335128, 24'd8022919, 24'd7783079, 24'd7663072, 24'd7686647, 24'd7849139, 24'd8118391, 24'd8441118, 24'd8753454, 24'd8993587, 24'd9113995, 24'd9090851, 24'd8928734, 24'd8659727, 24'd8337066, 24'd8024605, 24'd7784179, 24'd7663369, 24'd7686082, 24'd7847823, 24'd8116585, 24'd8439179, 
24'd8751766, 24'd8992484, 24'd9113696, 24'd9091414, 24'd8930048, 24'd8661533, 24'd8339005, 24'd8026294, 24'd7785284, 24'd7663671, 24'd7685521, 24'd7846511, 24'd8114781, 24'd8437240, 24'd8750075, 24'd8991377, 24'd9113391, 24'd9091972, 24'd8931359, 24'd8663336, 24'd8340944, 24'd8027986, 24'd7786393, 24'd7663978, 24'd7684965, 24'd7845202, 24'd8112978, 24'd8435301, 24'd8748383, 24'd8990266, 
24'd9113082, 24'd9092526, 24'd8932665, 24'd8665137, 24'd8342884, 24'd8029680, 24'd7787506, 24'd7664290, 24'd7684415, 24'd7843898, 24'd8111178, 24'd8433361, 24'd8746687, 24'd8989150, 24'd9112767, 24'd9093074, 24'd8933968, 24'd8666937, 24'd8344824, 24'd8031376, 24'd7788624, 24'd7664607, 24'd7683869, 24'd7842597, 24'd8109380, 24'd8431421, 24'd8744989, 24'd8988031, 24'd9112447, 24'd9093617, 
24'd8935267, 24'd8668734, 24'd8346764, 24'd8033075, 24'd7789746, 24'd7664930, 24'd7683328, 24'd7841300, 24'd8107583, 24'd8429480, 24'd8743289, 24'd8986907, 24'd9112122, 24'd9094156, 24'd8936562, 24'd8670529, 24'd8348705, 24'd8034777, 24'd7790872, 24'd7665257, 24'd7682792, 24'd7840007, 24'd8105789, 24'd8427540, 24'd8741586, 24'd8985779, 24'd9111792, 24'd9094689, 24'd8937853, 24'd8672323, 
24'd8350646, 24'd8036481, 24'd7792002, 24'd7665589, 24'd7682261, 24'd7838717, 24'd8103996, 24'd8425599, 24'd8739881, 24'd8984647, 24'd9111457, 24'd9095218, 24'd8939141, 24'd8674114, 24'd8352587, 24'd8038188, 24'd7793136, 24'd7665927, 24'd7681735, 24'd7837432, 24'd8102206, 24'd8423657, 24'd8738173, 24'd8983510, 24'd9111117, 24'd9095741, 24'd8940424, 24'd8675904, 24'd8354528, 24'd8039897, 
24'd7794274, 24'd7666270, 24'd7681214, 24'd7836150, 24'd8100417, 24'd8421716, 24'd8736463, 24'd8982370, 24'd9110772, 24'd9096260, 24'd8941704, 24'd8677692, 24'd8356470, 24'd8041608, 24'd7795417, 24'd7666617, 24'd7680698, 24'd7834873, 24'd8098631, 24'd8419774, 24'd8734750, 24'd8981225, 24'd9110422, 24'd9096773, 24'd8942980, 24'd8679477, 24'd8358412, 24'd8043322, 24'd7796564, 24'd7666970, 
24'd7680187, 24'd7833599, 24'd8096846, 24'd8417832, 24'd8733035, 24'd8980076, 24'd9110067, 24'd9097282, 24'd8944252, 24'd8681260, 24'd8360354, 24'd8045038, 24'd7797715, 24'd7667328, 24'd7679681, 24'd7832329, 24'd8095064, 24'd8415890, 24'd8731318, 24'd8978923, 24'd9109707, 24'd9097786, 24'd8945520, 24'd8683042, 24'd8362296, 24'd8046757, 24'd7798870, 24'd7667691, 24'd7679179, 24'd7831063, 
24'd8093283, 24'd8413948, 24'd8729598, 24'd8977766, 24'd9109341, 24'd9098284, 24'd8946784, 24'd8684821, 24'd8364238, 24'd8048478, 24'd7800029, 24'd7668058, 24'd7678683, 24'd7829801, 24'd8091505, 24'd8412005, 24'd8727875, 24'd8976605, 24'd9108971, 24'd9098778, 24'd8948044, 24'd8686598, 24'd8366181, 24'd8050202, 24'd7801192, 24'd7668431, 24'd7678192, 24'd7828542, 24'd8089729, 24'd8410063, 
24'd8726151, 24'd8975439, 24'd9108595, 24'd9099267, 24'd8949300, 24'd8688374, 24'd8368124, 24'd8051928, 24'd7802360, 24'd7668809, 24'd7677706, 24'd7827288, 24'd8087955, 24'd8408120, 24'd8724424, 24'd8974270, 24'd9108215, 24'd9099751, 24'd8950553, 24'd8690147, 24'd8370067, 24'd8053656, 24'd7803531, 24'd7669192, 24'd7677224, 24'd7826038, 24'd8086183, 24'd8406177, 24'd8722694, 24'd8973096, 
24'd9107829, 24'd9100229, 24'd8951801, 24'd8691918, 24'd8372010, 24'd8055386, 24'd7804707, 24'd7669580, 24'd7676748, 24'd7824791, 24'd8084413, 24'd8404234, 24'd8720962, 24'd8971919, 24'd9107439, 24'd9100703, 24'd8953045, 24'd8693686, 24'd8373953, 24'd8057119, 24'd7805887, 24'd7669974, 24'd7676277, 24'd7823549, 24'd8082645, 24'd8402291, 24'd8719228, 24'd8970737, 24'd9107043, 24'd9101172, 
24'd8954286, 24'd8695453, 24'd8375896, 24'd8058855, 24'd7807071, 24'd7670372, 24'd7675810, 24'd7822310, 24'd8080879, 24'd8400347, 24'd8717492, 24'd8969551, 24'd9106642, 24'd9101636, 24'd8955522, 24'd8697218, 24'd8377839, 24'd8060592, 24'd7808259, 24'd7670775, 24'd7675349, 24'd7821076, 24'd8079116, 24'd8398404, 24'd8715753, 24'd8968361, 24'd9106237, 24'd9102095, 24'd8956755, 24'd8698980, 
24'd8379783, 24'd8062332, 24'd7809451, 24'd7671183, 24'd7674893, 24'd7819845, 24'd8077355, 24'd8396461, 24'd8714012, 24'd8967167, 24'd9105826, 24'd9102548, 24'd8957983, 24'd8700740, 24'd8381726, 24'd8064074, 24'd7810647, 24'd7671596, 24'd7674442, 24'd7818619, 24'd8075596, 24'd8394517, 24'd8712269, 24'd8965969, 24'd9105410, 24'd9102997, 24'd8959208, 24'd8702498, 24'd8383670, 24'd8065819, 
24'd7811847, 24'd7672015, 24'd7673995, 24'd7817396, 24'd8073839, 24'd8392574, 24'd8710523, 24'd8964767, 24'd9104989, 24'd9103441, 24'd8960429, 24'd8704254, 24'd8385613, 24'd8067565, 24'd7813051, 24'd7672438, 24'd7673554, 24'd7816178, 24'd8072084, 24'd8390630, 24'd8708776, 24'd8963561, 24'd9104563, 24'd9103880, 24'd8961645, 24'd8706007, 24'd8387557, 24'd8069314, 24'd7814259, 24'd7672866, 
24'd7673118, 24'd7814963, 24'd8070332, 24'd8388686, 24'd8707026, 24'd8962350, 24'd9104133, 24'd9104314, 24'd8962858, 24'd8707759, 24'd8389500, 24'd8071065, 24'd7815471, 24'd7673300, 24'd7672686, 24'd7813753, 24'd8068581, 24'd8386743, 24'd8705273, 24'd8961136, 24'd9103697, 24'd9104742, 24'd8964066, 24'd8709508, 24'd8391444, 24'd8072819, 24'd7816687, 24'd7673738, 24'd7672260, 24'd7812546, 
24'd8066833, 24'd8384799, 24'd8703519, 24'd8959918, 24'd9103256, 24'd9105166, 24'd8965271, 24'd8711255, 24'd8393387, 24'd8074574, 24'd7817908, 24'd7674182, 24'd7671839, 24'd7811344, 24'd8065088, 24'd8382856, 24'd8701762, 24'd8958696, 24'd9102810, 24'd9105585, 24'd8966471, 24'd8712999, 24'd8395331, 24'd8076332, 24'd7819132, 24'd7674630, 24'd7671423, 24'd7810145, 24'd8063344, 24'd8380912, 
24'd8700003, 24'd8957469, 24'd9102359, 24'd9105998, 24'd8967667, 24'd8714742, 24'd8397274, 24'd8078092, 24'd7820360, 24'd7675083, 24'd7671012, 24'd7808951, 24'd8061603, 24'd8378969, 24'd8698242, 24'd8956239, 24'd9101903, 24'd9106407, 24'd8968860, 24'd8716482, 24'd8399218, 24'd8079854, 24'd7821592, 24'd7675542, 24'd7670606, 24'd7807761, 24'd8059864, 24'd8377025, 24'd8696479, 24'd8955005, 
24'd9101442, 24'd9106811, 24'd8970048, 24'd8718219, 24'd8401161, 24'd8081619, 24'd7822829, 24'd7676005, 24'd7670204, 24'd7806574, 24'd8058128, 24'd8375082, 24'd8694713, 24'd8953767, 24'd9100976, 24'd9107209, 24'd8971232, 24'd8719955, 24'd8403104, 24'd8083385, 24'd7824069, 24'd7676474, 24'd7669808, 24'd7805392, 24'd8056393, 24'd8373139, 24'd8692946, 24'd8952525, 24'd9100505, 24'd9107603, 
24'd8972412, 24'd8721688, 24'd8405048, 24'd8085154, 24'd7825313, 24'd7676947, 24'd7669417, 24'd7804214, 24'd8054661, 24'd8371196, 24'd8691176, 24'd8951279, 24'd9100029, 24'd9107991, 24'd8973588, 24'd8723419, 24'd8406991, 24'd8086925, 24'd7826561, 24'd7677425, 24'd7669031, 24'd7803040, 24'd8052932, 24'd8369253, 24'd8689404, 24'd8950029, 24'd9099549, 24'd9108375, 24'd8974760, 24'd8725147, 
24'd8408934, 24'd8088697, 24'd7827813, 24'd7677909, 24'd7668650, 24'd7801870, 24'd8051204, 24'd8367310, 24'd8687630, 24'd8948775, 24'd9099063, 24'd9108753, 24'd8975928, 24'd8726873, 24'd8410876, 24'd8090472, 24'd7829069, 24'd7678397, 24'd7668275, 24'd7800705, 24'd8049480, 24'd8365367, 24'd8685854, 24'd8947517, 24'd9098572, 24'd9109126, 24'd8977092, 24'd8728597, 24'd8412819, 24'd8092249, 
24'd7830329, 24'd7678890, 24'd7667904, 24'd7799543, 24'd8047757, 24'd8363425, 24'd8684076, 24'd8946255, 24'd9098076, 24'd9109495, 24'd8978251, 24'd8730318, 24'd8414761, 24'd8094029, 24'd7831593, 24'd7679389, 24'd7667538, 24'd7798386, 24'd8046037, 24'd8361483, 24'd8682296, 24'd8944989, 24'd9097575, 24'd9109858, 24'd8979407, 24'd8732037, 24'd8416704, 24'd8095810, 24'd7832860, 24'd7679892, 
24'd7667177, 24'd7797232, 24'd8044319, 24'd8359540, 24'd8680514, 24'd8943719, 24'd9097070, 24'd9110216, 24'd8980558, 24'd8733754, 24'd8418646, 24'd8097593, 24'd7834132, 24'd7680400, 24'd7666822, 24'd7796083, 24'd8042604, 24'd8357598, 24'd8678729, 24'd8942446, 24'd9096559, 24'd9110569, 24'd8981705, 24'd8735468, 24'd8420587, 24'd8099378, 24'd7835407, 24'd7680913, 24'd7666471, 24'd7794938, 
24'd8040891, 24'd8355657, 24'd8676943, 24'd8941169, 24'd9096043, 24'd9110917, 24'd8982848, 24'd8737179, 24'd8422529, 24'd8101166, 24'd7836687, 24'd7681432, 24'd7666125, 24'd7793797, 24'd8039181, 24'd8353715, 24'd8675155, 24'd8939887, 24'd9095522, 24'd9111260, 24'd8983987, 24'd8738889, 24'd8424470, 24'd8102955, 24'd7837970, 24'd7681955, 24'd7665785, 24'd7792660, 24'd8037473, 24'd8351774, 
24'd8673364, 24'd8938602, 24'd9094997, 24'd9111598, 24'd8985121, 24'd8740595, 24'd8426412, 24'd8104746, 24'd7839257, 24'd7682483, 24'd7665450, 24'd7791528, 24'd8035767, 24'd8349833, 24'd8671572, 24'd8937313, 24'd9094466, 24'd9111931, 24'd8986252, 24'd8742300, 24'd8428352, 24'd8106540, 24'd7840548, 24'd7683016, 24'd7665119, 24'd7790400, 24'd8034064, 24'd8347892, 24'd8669778, 24'd8936020, 
24'd9093931, 24'd9112259, 24'd8987378, 24'd8744001, 24'd8430293, 24'd8108335, 24'd7841843, 24'd7683554, 24'd7664794, 24'd7789275, 24'd8032364, 24'd8345952, 24'd8667981, 24'd8934724, 24'd9093390, 24'd9112582, 24'd8988500, 24'd8745701, 24'd8432233, 24'd8110132, 24'd7843141, 24'd7684097, 24'd7664474, 24'd7788155, 24'd8030665, 24'd8344012, 24'd8666183, 24'd8933423, 24'd9092845, 24'd9112899, 
24'd8989618, 24'd8747398, 24'd8434173, 24'd8111932, 24'd7844444, 24'd7684645, 24'd7664159, 24'd7787040, 24'd8028970, 24'd8342072, 24'd8664383, 24'd8932119, 24'd9092295, 24'd9113212, 24'd8990732, 24'd8749092, 24'd8436113, 24'd8113733, 24'd7845750, 24'd7685197, 24'd7663849, 24'd7785928, 24'd8027277, 24'd8340132, 24'd8662581, 24'd8930811, 24'd9091739, 24'd9113520, 24'd8991841, 24'd8750784, 
24'd8438052, 24'd8115536, 24'd7847060, 24'd7685755, 24'd7663544, 24'd7784821, 24'd8025586, 24'd8338193, 24'd8660777, 24'd8929499, 24'd9091179, 24'd9113822, 24'd8992946, 24'd8752473, 24'd8439991, 24'd8117341, 24'd7848374, 24'd7686318, 24'd7663244, 24'd7783718, 24'd8023898, 24'd8336254, 24'd8658971, 24'd8928183, 24'd9090614, 24'd9114119, 24'd8994047, 24'd8754160, 24'd8441930, 24'd8119148, 
24'd7849691, 24'd7686885, 24'd7662949, 24'd7782619, 24'd8022213, 24'd8334316, 24'd8657163, 24'd8926863, 24'd9090044, 24'd9114411, 24'd8995144, 24'd8755844, 24'd8443868, 24'd8120957, 24'd7851013, 24'd7687458, 24'd7662659, 24'd7781524, 24'd8020530, 24'd8332378, 24'd8655353, 24'd8925540, 24'd9089469, 24'd9114699, 24'd8996236, 24'd8757525, 24'd8445806, 24'd8122767, 24'd7852338, 24'd7688035, 
24'd7662375, 24'd7780434, 24'd8018850, 24'd8330440, 24'd8653542, 24'd8924213, 24'd9088889, 24'd9114981, 24'd8997324, 24'd8759204, 24'd8447744, 24'd8124580, 24'd7853667, 24'd7688618, 24'd7662095, 24'd7779348, 24'd8017172, 24'd8328503, 24'd8651728, 24'd8922882, 24'd9088304, 24'd9115258, 24'd8998408, 24'd8760881, 24'd8449681, 24'd8126394, 24'd7855000, 24'd7689205, 24'd7661821, 24'd7778266, 
24'd8015497, 24'd8326566, 24'd8649913, 24'd8921548, 24'd9087715, 24'd9115530, 24'd8999488, 24'd8762554, 24'd8451617, 24'd8128211, 24'd7856336, 24'd7689797, 24'd7661551, 24'd7777189, 24'd8013825, 24'd8324630, 24'd8648096, 24'd8920209, 24'd9087120, 24'd9115796, 24'd9000563, 24'd8764225, 24'd8453553, 24'd8130029, 24'd7857676, 24'd7690394, 24'd7661287, 24'd7776116, 24'd8012155, 24'd8322694, 
24'd8646277, 24'd8918867, 24'd9086520, 24'd9116058, 24'd9001634, 24'd8765894, 24'd8455489, 24'd8131849, 24'd7859020, 24'd7690996, 24'd7661028, 24'd7775047, 24'd8010488, 24'd8320758, 24'd8644456, 24'd8917521, 24'd9085916, 24'd9116315, 24'd9002701, 24'd8767560, 24'd8457424, 24'd8133670, 24'd7860368, 24'd7691603, 24'd7660774, 24'd7773982, 24'd8008823, 24'd8318823, 24'd8642633, 24'd8916172, 
24'd9085307, 24'd9116566, 24'd9003764, 24'd8769223, 24'd8459359, 24'd8135494, 24'd7861719, 24'd7692215, 24'd7660525, 24'd7772922, 24'd8007161, 24'd8316889, 24'd8640809, 24'd8914819, 24'd9084693, 24'd9116812, 24'd9004822, 24'd8770883, 24'd8461293, 24'd8137319, 24'd7863074, 24'd7692831, 24'd7660281, 24'd7771866, 24'd8005502, 24'd8314955, 24'd8638983, 24'd8913462, 24'd9084074, 24'd9117054, 
24'd9005876, 24'd8772541, 24'd8463227, 24'd8139146, 24'd7864433, 24'd7693453, 24'd7660043, 24'd7770814, 24'd8003846, 24'd8313021, 24'd8637155, 24'd8912101, 24'd9083450, 24'd9117290, 24'd9006925, 24'd8774196, 24'd8465160, 24'd8140975, 24'd7865795, 24'd7694079, 24'd7659809, 24'd7769767, 24'd8002192, 24'd8311088, 24'd8635325, 24'd8910737, 24'd9082821, 24'd9117521, 24'd9007970, 24'd8775849, 
24'd8467093, 24'd8142805, 24'd7867161, 24'd7694710, 24'd7659581, 24'd7768724, 24'd8000541, 24'd8309156, 24'd8633494, 24'd8909369, 24'd9082187, 24'd9117747, 24'd9009011, 24'd8777499, 24'd8469025, 24'd8144637, 24'd7868531, 24'd7695346, 24'd7659357, 24'd7767685, 24'd7998893, 24'd8307224, 24'd8631661, 24'd8907998, 24'd9081549, 24'd9117968, 24'd9010048, 24'd8779146, 24'd8470957, 24'd8146471, 
24'd7869904, 24'd7695987, 24'd7659139, 24'd7766651, 24'd7997247, 24'd8305293, 24'd8629826, 24'd8906623, 24'd9080905, 24'd9118183, 24'd9011080, 24'd8780790, 24'd8472888, 24'd8148307, 24'd7871281, 24'd7696633, 24'd7658926, 24'd7765621, 24'd7995604, 24'd8303362, 24'd8627990, 24'd8905244, 24'd9080257, 24'd9118394, 24'd9012107, 24'd8782431, 24'd8474818, 24'd8150144, 24'd7872662, 24'd7697284, 
24'd7658718, 24'd7764595, 24'd7993964, 24'd8301432, 24'd8626151, 24'd8903862, 24'd9079604, 24'd9118599, 24'd9013131, 24'd8784070, 24'd8476748, 24'd8151983, 24'd7874046, 24'd7697939, 24'd7658515, 24'd7763574, 24'd7992327, 24'd8299502, 24'd8624312, 24'd8902476, 24'd9078946, 24'd9118800, 24'd9014150, 24'd8785706, 24'd8478677, 24'd8153824, 24'd7875434, 24'd7698600, 24'd7658317, 24'd7762557, 
24'd7990692, 24'd8297573, 24'd8622470, 24'd8901086, 24'd9078283, 24'd9118995, 24'd9015164, 24'd8787339, 24'd8480606, 24'd8155666, 24'd7876825, 24'd7699265, 24'd7658124, 24'd7761545, 24'd7989060, 24'd8295645, 24'd8620627, 24'd8899693, 24'd9077616, 24'd9119185, 24'd9016175, 24'd8788970, 24'd8482534, 24'd8157510, 24'd7878220, 24'd7699935, 24'd7657937, 24'd7760537, 24'd7987431, 24'd8293717, 
24'd8618782, 24'd8898296, 24'd9076943, 24'd9119370, 24'd9017180, 24'd8790597, 24'd8484461, 24'd8159356, 24'd7879619, 24'd7700610, 24'd7657754, 24'd7759533, 24'd7985805, 24'd8291790, 24'd8616936, 24'd8896896, 24'd9076266, 24'd9119550, 24'd9018182, 24'd8792222, 24'd8486388, 24'd8161203, 24'd7881021, 24'd7701290, 24'd7657577, 24'd7758534, 24'd7984182, 24'd8289864, 24'd8615088, 24'd8895492, 
24'd9075584, 24'd9119725, 24'd9019179, 24'd8793844, 24'd8488314, 24'd8163052, 24'd7882427, 24'd7701974, 24'd7657405, 24'd7757539, 24'd7982561, 24'd8287939, 24'd8613238, 24'd8894084, 24'd9074897, 24'd9119894, 24'd9020171, 24'd8795463, 24'd8490239, 24'd8164902, 24'd7883836, 24'd7702663, 24'd7657238, 24'd7756549, 24'd7980943, 24'd8286014, 24'd8611387, 24'd8892673, 24'd9074205, 24'd9120059, 
24'd9021160, 24'd8797079, 24'd8492163, 24'd8166754, 24'd7885249, 24'd7703357, 24'd7657076, 24'd7755563, 24'd7979329, 24'd8284090, 24'd8609535, 24'd8891259, 24'd9073509, 24'd9120218, 24'd9022143, 24'd8798693, 24'd8494087, 24'd8168607, 24'd7886665, 24'd7704056, 24'd7656919, 24'd7754582, 24'd7977717, 24'd8282166, 24'd8607680, 24'd8889840, 24'd9072807, 24'd9120372, 24'd9023123, 24'd8800303, 
24'd8496010, 24'd8170462, 24'd7888085, 24'd7704760, 24'd7656767, 24'd7753605, 24'd7976108, 24'd8280244, 24'd8605825, 24'd8888419, 24'd9072101, 24'd9120522, 24'd9024097, 24'd8801911, 24'd8497932, 24'd8172319, 24'd7889508, 24'd7705469, 24'd7656621, 24'd7752632, 24'd7974501, 24'd8278322, 24'd8603967, 24'd8886994, 24'd9071390, 24'd9120665, 24'd9025068, 24'd8803516, 24'd8499854, 24'd8174177, 
24'd7890935, 24'd7706182, 24'd7656479, 24'd7751664, 24'd7972898, 24'd8276401, 24'd8602109, 24'd8885565, 24'd9070675, 24'd9120804, 24'd9026034, 24'd8805117, 24'd8501775, 24'd8176036, 24'd7892365, 24'd7706900, 24'd7656343, 24'd7750700, 24'd7971298, 24'd8274480, 24'd8600248, 24'd8884133, 24'd9069954, 24'd9120938, 24'd9026995, 24'd8806716, 24'd8503695, 24'd8177897, 24'd7893799, 24'd7707623, 
24'd7656212, 24'd7749741, 24'd7969700, 24'd8272561, 24'd8598387, 24'd8882697, 24'd9069229, 24'd9121067, 24'd9027952, 24'd8808312, 24'd8505614, 24'd8179760, 24'd7895237, 24'd7708351, 24'd7656086, 24'd7748786, 24'd7968106, 24'd8270642, 24'd8596523, 24'd8881258, 24'd9068499, 24'd9121190, 24'd9028904, 24'd8809905, 24'd8507532, 24'd8181624, 24'd7896677, 24'd7709083, 24'd7655965, 24'd7747836, 
24'd7966514, 24'd8268724, 24'd8594659, 24'd8879816, 24'd9067764, 24'd9121308, 24'd9029852, 24'd8811495, 24'd8509450, 24'd8183489, 24'd7898122, 24'd7709820, 24'd7655849, 24'd7746890, 24'd7964926, 24'd8266807, 24'd8592792, 24'd8878370, 24'd9067024, 24'd9121421, 24'd9030796, 24'd8813082, 24'd8511366, 24'd8185356, 24'd7899569, 24'd7710562, 24'd7655739, 24'd7745949, 24'd7963340, 24'd8264891, 
24'd8590925, 24'd8876921, 24'd9066280, 24'd9121530, 24'd9031735, 24'd8814667, 24'd8513282, 24'd8187224, 24'd7901020, 24'd7711309, 24'd7655633, 24'd7745012, 24'd7961757, 24'd8262976, 24'd8589056, 24'd8875468, 24'd9065531, 24'd9121632, 24'd9032669, 24'd8816248, 24'd8515197, 24'd8189094, 24'd7902475, 24'd7712060, 24'd7655533, 24'd7744080, 24'd7960178, 24'd8261061, 24'd8587185, 24'd8874012, 
24'd9064777, 24'd9121730, 24'd9033599, 24'd8817826, 24'd8517111, 24'd8190965, 24'd7903933, 24'd7712816, 24'd7655438, 24'd7743152, 24'd7958601, 24'd8259147, 24'd8585314, 24'd8872552, 24'd9064019, 24'd9121823, 24'd9034525, 24'd8819401, 24'd8519024, 24'd8192838, 24'd7905394, 24'd7713577, 24'd7655348, 24'd7742229, 24'd7957028, 24'd8257235, 24'd8583441, 24'd8871089, 24'd9063255, 24'd9121910, 
24'd9035446, 24'd8820973, 24'd8520936, 24'd8194712, 24'd7906859, 24'd7714343, 24'd7655263, 24'd7741311, 24'd7955457, 24'd8255323, 24'd8581566, 24'd8869623, 24'd9062487, 24'd9121993, 24'd9036362, 24'd8822542, 24'd8522847, 24'd8196587, 24'd7908327, 24'd7715113, 24'd7655183, 24'd7740396, 24'd7953889, 24'd8253412, 24'd8579690, 24'd8868153, 24'd9061715, 24'd9122070, 24'd9037274, 24'd8824108, 
24'd8524758, 24'd8198463, 24'd7909798, 24'd7715888, 24'd7655109, 24'd7739487, 24'd7952325, 24'd8251502, 24'd8577813, 24'd8866680, 24'd9060937, 24'd9122142, 24'd9038181, 24'd8825671, 24'd8526667, 24'd8200341, 24'd7911273, 24'd7716668, 24'd7655039, 24'd7738582, 24'd7950763, 24'd8249594, 24'd8575934, 24'd8865203, 24'd9060155, 24'd9122209, 24'd9039084, 24'd8827231, 24'd8528576, 24'd8202220, 
24'd7912751, 24'd7717453, 24'd7654975, 24'd7737681, 24'd7949205, 24'd8247686, 24'd8574054, 24'd8863724, 24'd9059368, 24'd9122270, 24'd9039982, 24'd8828788, 24'd8530483, 24'd8204101, 24'd7914233, 24'd7718242, 24'd7654916, 24'd7736786, 24'd7947650, 24'd8245779, 24'd8572173, 24'd8862240, 24'd9058577, 24'd9122327, 24'd9040876, 24'd8830342, 24'd8532389, 24'd8205983, 24'd7915717, 24'd7719036, 
24'd7654862, 24'd7735894, 24'd7946098, 24'd8243873, 24'd8570291, 24'd8860754, 24'd9057780, 24'd9122378, 24'd9041765, 24'd8831892, 24'd8534295, 24'd8207866, 24'd7917205, 24'd7719835, 24'd7654813, 24'd7735007, 24'd7944548, 24'd8241968, 24'd8568407, 24'd8859264, 24'd9056979, 24'd9122425, 24'd9042649, 24'd8833440, 24'd8536199, 24'd8209750, 24'd7918697, 24'd7720638, 24'd7654769, 24'd7734125, 
24'd7943002, 24'd8240064, 24'd8566522, 24'd8857771, 24'd9056174, 24'd9122466, 24'd9043529, 24'd8834984, 24'd8538103, 24'd8211636, 24'd7920192, 24'd7721446, 24'd7654730, 24'd7733248, 24'd7941460, 24'd8238161, 24'd8564636, 24'd8856275, 24'd9055363, 24'd9122502, 24'd9044404, 24'd8836526, 24'd8540005, 24'd8213523, 24'd7921690, 24'd7722259, 24'd7654697, 24'd7732375, 24'd7939920, 24'd8236259, 
24'd8562748, 24'd8854775, 24'd9054548, 24'd9122533, 24'd9045275, 24'd8838064, 24'd8541906, 24'd8215411, 24'd7923191, 24'd7723076, 24'd7654669, 24'd7731506, 24'd7938383, 24'd8234359, 24'd8560860, 24'd8853272, 24'd9053729, 24'd9122559, 24'd9046141, 24'd8839599, 24'd8543806, 24'd8217300, 24'd7924695, 24'd7723898, 24'd7654645, 24'd7730643, 24'd7936850, 24'd8232459, 24'd8558970, 24'd8851766, 
24'd9052904, 24'd9122579, 24'd9047003, 24'd8841131, 24'd8545705, 24'd8219191, 24'd7926203, 24'd7724725, 24'd7654627, 24'd7729783, 24'd7935320, 24'd8230561, 24'd8557079, 24'd8850257, 24'd9052075, 24'd9122595, 24'd9047859, 24'd8842659, 24'd8547603, 24'd8221082, 24'd7927714, 24'd7725556, 24'd7654615, 24'd7728929, 24'd7933792, 24'd8228663, 24'd8555186, 24'd8848744, 24'd9051241, 24'd9122605, 
24'd9048712, 24'd8844185, 24'd8549500, 24'd8222975, 24'd7929229, 24'd7726392, 24'd7654607, 24'd7728079, 24'd7932269, 24'd8226767, 24'd8553293, 24'd8847228, 24'd9050403, 24'd9122610, 24'd9049559, 24'd8845707, 24'd8551396, 24'd8224869, 24'd7930746, 24'd7727233, 24'd7654604, 24'd7727234, 24'd7930748, 24'd8224872, 24'd8551398, 24'd8845709, 24'd9049560, 24'd9122610, 24'd9050402, 24'd8847226, 
24'd8553291, 24'd8226764, 24'd7932267, 24'd7728078, 24'd7654607, 24'd7726393, 24'd7929230, 24'd8222978, 24'd8549503, 24'd8844187, 24'd9048713, 24'd9122605, 24'd9051240, 24'd8848742, 24'd8555184, 24'd8228661, 24'd7933791, 24'd7728928, 24'd7654615, 24'd7725557, 24'd7927716, 24'd8221085, 24'd8547606, 24'd8842661, 24'd9047860, 24'd9122595, 24'd9052074, 24'd8850255, 24'd8557076, 24'd8230558, 
24'd7935318, 24'd7729782, 24'd7654627, 24'd7724726, 24'd7926205, 24'd8219193, 24'd8545708, 24'd8841133, 24'd9047004, 24'd9122579, 24'd9052903, 24'd8851764, 24'd8558967, 24'd8232457, 24'd7936848, 24'd7730642, 24'd7654645, 24'd7723899, 24'd7924697, 24'd8217303, 24'd8543809, 24'd8839601, 24'd9046142, 24'd9122559, 24'd9053727, 24'd8853270, 24'd8560857, 24'd8234356, 24'd7938381, 24'd7731505, 
24'd7654669, 24'd7723077, 24'd7923193, 24'd8215413, 24'd8541908, 24'd8838066, 24'd9045276, 24'd9122533, 24'd9054547, 24'd8854773, 24'd8562746, 24'd8236257, 24'd7939918, 24'd7732374, 24'd7654697, 24'd7722260, 24'd7921692, 24'd8213525, 24'd8540007, 24'd8836528, 24'd9044405, 24'd9122502, 24'd9055362, 24'd8856273, 24'd8564633, 24'd8238159, 24'd7941458, 24'd7733247, 24'd7654730, 24'd7721447, 
24'd7920193, 24'd8211638, 24'd8538105, 24'd8834986, 24'd9043530, 24'd9122466, 24'd9056173, 24'd8857769, 24'd8566520, 24'd8240062, 24'd7943001, 24'd7734124, 24'd7654769, 24'd7720639, 24'd7918699, 24'd8209753, 24'd8536202, 24'd8833442, 24'd9042650, 24'd9122425, 24'd9056978, 24'd8859262, 24'd8568405, 24'd8241966, 24'd7944547, 24'd7735006, 24'd7654813, 24'd7719836, 24'd7917207, 24'd8207868, 
24'd8534297, 24'd8831894, 24'd9041766, 24'd9122379, 24'd9057779, 24'd8860752, 24'd8570288, 24'd8243870, 24'd7946096, 24'd7735893, 24'd7654862, 24'd7719037, 24'd7915719, 24'd8205985, 24'd8532392, 24'd8830344, 24'd9040877, 24'd9122327, 24'd9058576, 24'd8862239, 24'd8572171, 24'd8245776, 24'd7947648, 24'd7736784, 24'd7654916, 24'd7718243, 24'd7914234, 24'd8204103, 24'd8530485, 24'd8828790, 
24'd9039983, 24'd9122270, 24'd9059367, 24'd8863722, 24'd8574052, 24'd8247683, 24'd7949203, 24'd7737680, 24'd7654975, 24'd7717454, 24'd7912753, 24'd8202223, 24'd8528578, 24'd8827233, 24'd9039085, 24'd9122209, 24'd9060154, 24'd8865202, 24'd8575932, 24'd8249591, 24'd7950761, 24'd7738581, 24'd7655039, 24'd7716669, 24'd7911275, 24'd8200344, 24'd8526669, 24'd8825673, 24'd9038182, 24'd9122142, 
24'd9060936, 24'd8866678, 24'd8577810, 24'd8251500, 24'd7952323, 24'd7739486, 24'd7655109, 24'd7715889, 24'd7909800, 24'd8198466, 24'd8524760, 24'd8824110, 24'd9037275, 24'd9122070, 24'd9061714, 24'd8868151, 24'd8579688, 24'd8253410, 24'd7953887, 24'd7740395, 24'd7655183, 24'd7715114, 24'd7908329, 24'd8196589, 24'd8522850, 24'd8822544, 24'd9036363, 24'd9121993, 24'd9062486, 24'd8869621, 
24'd8581564, 24'd8255321, 24'd7955455, 24'd7741309, 24'd7655263, 24'd7714344, 24'd7906861, 24'd8194714, 24'd8520939, 24'd8820975, 24'd9035447, 24'd9121910, 24'd9063254, 24'd8871087, 24'd8583438, 24'd8257232, 24'd7957026, 24'd7742228, 24'd7655348, 24'd7713578, 24'd7905396, 24'd8192840, 24'd8519026, 24'd8819403, 24'd9034526, 24'd9121823, 24'd9064018, 24'd8872550, 24'd8585311, 24'd8259145, 
24'd7958599, 24'd7743151, 24'd7655438, 24'd7712817, 24'd7903935, 24'd8190968, 24'd8517113, 24'd8817828, 24'd9033601, 24'd9121730, 24'd9064776, 24'd8874010, 24'd8587183, 24'd8261059, 24'd7960176, 24'd7744079, 24'd7655533, 24'd7712061, 24'd7902477, 24'd8189096, 24'd8515199, 24'd8816250, 24'd9032671, 24'd9121633, 24'd9065530, 24'd8875466, 24'd8589054, 24'd8262973, 24'd7961755, 24'd7745011, 
24'd7655633, 24'd7711310, 24'd7901022, 24'd8187227, 24'd8513284, 24'd8814669, 24'd9031736, 24'd9121530, 24'd9066279, 24'd8876919, 24'd8590923, 24'd8264888, 24'd7963338, 24'd7745948, 24'd7655739, 24'd7710563, 24'd7899571, 24'd8185359, 24'd8511369, 24'd8813084, 24'd9030797, 24'd9121422, 24'd9067024, 24'd8878368, 24'd8592790, 24'd8266805, 24'd7964924, 24'd7746889, 24'd7655849, 24'd7709821, 
24'd7898123, 24'd8183492, 24'd8509452, 24'd8811497, 24'd9029854, 24'd9121308, 24'd9067763, 24'd8879814, 24'd8594656, 24'd8268722, 24'd7966512, 24'd7747835, 24'd7655965, 24'd7709084, 24'd7896679, 24'd8181626, 24'd8507534, 24'd8809907, 24'd9028906, 24'd9121190, 24'd9068498, 24'd8881257, 24'd8596521, 24'd8270640, 24'd7968104, 24'd7748785, 24'd7656086, 24'd7708351, 24'd7895238, 24'd8179762, 
24'd8505616, 24'd8808314, 24'd9027953, 24'd9121067, 24'd9069228, 24'd8882696, 24'd8598384, 24'd8272558, 24'd7969698, 24'd7749740, 24'd7656212, 24'd7707624, 24'd7893801, 24'd8177900, 24'd8503697, 24'd8806718, 24'd9026996, 24'd9120938, 24'd9069953, 24'd8884131, 24'd8600246, 24'd8274478, 24'd7971296, 24'd7750699, 24'd7656343, 24'd7706901, 24'd7892367, 24'd8176039, 24'd8501777, 24'd8805119, 
24'd9026035, 24'd9120804, 24'd9070674, 24'd8885563, 24'd8602106, 24'd8276398, 24'd7972896, 24'd7751663, 24'd7656479, 24'd7706183, 24'd7890937, 24'd8174179, 24'd8499856, 24'd8803518, 24'd9025069, 24'd9120666, 24'd9071389, 24'd8886992, 24'd8603965, 24'd8278319, 24'd7974499, 24'd7752631, 24'd7656621, 24'd7705470, 24'd7889510, 24'd8172321, 24'd8497935, 24'd8801913, 24'd9024099, 24'd9120522, 
24'd9072100, 24'd8888417, 24'd8605822, 24'd8280241, 24'd7976106, 24'd7753603, 24'd7656767, 24'd7704761, 24'd7888087, 24'd8170465, 24'd8496013, 24'd8800305, 24'd9023124, 24'd9120373, 24'd9072806, 24'd8889839, 24'd8607678, 24'd8282164, 24'd7977715, 24'd7754580, 24'd7656919, 24'd7704057, 24'd7886667, 24'd8168610, 24'd8494090, 24'd8798695, 24'd9022144, 24'd9120218, 24'd9073508, 24'd8891257, 
24'd8609532, 24'd8284087, 24'd7979327, 24'd7755562, 24'd7657076, 24'd7703358, 24'd7885251, 24'd8166756, 24'd8492166, 24'd8797081, 24'd9021161, 24'd9120059, 24'd9074204, 24'd8892671, 24'd8611385, 24'd8286011, 24'd7980941, 24'd7756548, 24'd7657238, 24'd7702664, 24'd7883838, 24'd8164904, 24'd8490241, 24'd8795465, 24'd9020173, 24'd9119895, 24'd9074896, 24'd8894082, 24'd8613236, 24'd8287936, 
24'd7982559, 24'd7757538, 24'd7657405, 24'd7701975, 24'd7882428, 24'd8163054, 24'd8488316, 24'd8793846, 24'd9019180, 24'd9119725, 24'd9075583, 24'd8895490, 24'd8615086, 24'd8289862, 24'd7984180, 24'd7758533, 24'd7657577, 24'd7701290, 24'd7881023, 24'd8161205, 24'd8486390, 24'd8792224, 24'd9018183, 24'd9119550, 24'd9076265, 24'd8896894, 24'd8616934, 24'd8291788, 24'd7985803, 24'd7759532, 
24'd7657754, 24'd7700611, 24'd7879621, 24'd8159358, 24'd8484464, 24'd8790599, 24'd9017182, 24'd9119370, 24'd9076942, 24'd8898294, 24'd8618780, 24'd8293715, 24'd7987429, 24'd7760536, 24'd7657937, 24'd7699936, 24'd7878222, 24'd8157512, 24'd8482536, 24'd8788972, 24'd9016176, 24'd9119185, 24'd9077615, 24'd8899691, 24'd8620625, 24'd8295643, 24'd7989058, 24'd7761544, 24'd7658124, 24'd7699266, 
24'd7876827, 24'd8155669, 24'd8480608, 24'd8787341, 24'd9015166, 24'd9118995, 24'd9078282, 24'd8901084, 24'd8622468, 24'd8297571, 24'd7990690, 24'd7762556, 24'd7658317, 24'd7698601, 24'd7875436, 24'd8153826, 24'd8478680, 24'd8785708, 24'd9014151, 24'd9118800, 24'd9078945, 24'd8902474, 24'd8624309, 24'd8299500, 24'd7992324, 24'd7763573, 24'd7658515, 24'd7697940, 24'd7874048, 24'd8151986, 
24'd8476751, 24'd8784072, 24'd9013132, 24'd9118600, 24'd9079603, 24'd8903860, 24'd8626149, 24'd8301429, 24'd7993962, 24'd7764594, 24'd7658717, 24'd7697285, 24'd7872664, 24'd8150147, 24'd8474821, 24'd8782433, 24'd9012109, 24'd9118394, 24'd9080256, 24'd8905242, 24'd8627987, 24'd8303359, 24'd7995602, 24'd7765620, 24'd7658925, 24'd7696634, 24'd7871283, 24'd8148309, 24'd8472890, 24'd8780792, 
24'd9011081, 24'd9118184, 24'd9080904, 24'd8906621, 24'd8629824, 24'd8305290, 24'd7997245, 24'd7766650, 24'd7659139, 24'd7695988, 24'd7869906, 24'd8146474, 24'd8470959, 24'd8779148, 24'd9010049, 24'd9117968, 24'd9081548, 24'd8907996, 24'd8631658, 24'd8307221, 24'd7998890, 24'd7767684, 24'd7659357, 24'd7695347, 24'd7868533, 24'd8144640, 24'd8469028, 24'd8777501, 24'd9009012, 24'd9117747, 
24'd9082186, 24'd8909368, 24'd8633492, 24'd8309153, 24'd8000539, 24'd7768723, 24'd7659580, 24'd7694711, 24'd7867163, 24'd8142808, 24'd8467096, 24'd8775851, 24'd9007972, 24'd9117521, 24'd9082820, 24'd8910736, 24'd8635323, 24'd8311086, 24'd8002190, 24'd7769765, 24'd7659809, 24'd7694080, 24'd7865797, 24'd8140977, 24'd8465163, 24'd8774199, 24'd9006926, 24'd9117290, 24'd9083449, 24'd8912100, 
24'd8637153, 24'd8313019, 24'd8003844, 24'd7770813, 24'd7660042, 24'd7693454, 24'd7864435, 24'd8139148, 24'd8463230, 24'd8772543, 24'd9005877, 24'd9117054, 24'd9084073, 24'd8913460, 24'd8638980, 24'd8314952, 24'd8005500, 24'd7771864, 24'd7660281, 24'd7692832, 24'd7863076, 24'd8137321, 24'd8461296, 24'd8770886, 24'd9004823, 24'd9116813, 24'd9084692, 24'd8914817, 24'd8640807, 24'd8316886, 
24'd8007159, 24'd7772920, 24'd7660525, 24'd7692215, 24'd7861721, 24'd8135496, 24'd8459362, 24'd8769225, 24'd9003765, 24'd9116566, 24'd9085306, 24'd8916170, 24'd8642631, 24'd8318821, 24'd8008821, 24'd7773981, 24'd7660774, 24'd7691604, 24'd7860369, 24'd8133673, 24'd8457427, 24'd8767562, 24'd9002702, 24'd9116315, 24'd9085915, 24'd8917520, 24'd8644453, 24'd8320756, 24'd8010486, 24'd7775045, 
24'd7661028, 24'd7690997, 24'd7859022, 24'd8131851, 24'd8455492, 24'd8765896, 24'd9001636, 24'd9116058, 24'd9086520, 24'd8918866, 24'd8646274, 24'd8322691, 24'd8012153, 24'd7776114, 24'd7661287, 24'd7690395, 24'd7857678, 24'd8130031, 24'd8453556, 24'd8764228, 24'd9000565, 24'd9115797, 24'd9087119, 24'd8920208, 24'd8648093, 24'd8324627, 24'd8013823, 24'd7777187, 24'd7661551, 24'd7689798, 
24'd7856338, 24'd8128213, 24'd8451620, 24'd8762556, 24'd8999489, 24'd9115530, 24'd9087714, 24'd8921546, 24'd8649910, 24'd8326564, 24'd8015495, 24'd7778265, 24'd7661820, 24'd7689206, 24'd7855001, 24'd8126397, 24'd8449683, 24'd8760883, 24'd8998410, 24'd9115258, 24'd9088304, 24'd8922880, 24'd8651726, 24'd8328500, 24'd8017170, 24'd7779347, 24'd7662095, 24'd7688618, 24'd7853669, 24'd8124582, 
24'd8447746, 24'd8759206, 24'd8997326, 24'd9114981, 24'd9088888, 24'd8924211, 24'd8653539, 24'd8330438, 24'd8018848, 24'd7780433, 24'd7662374, 24'd7688036, 24'd7852340, 24'd8122770, 24'd8445809, 24'd8757527, 24'd8996238, 24'd9114699, 24'd9089468, 24'd8925538, 24'd8655351, 24'd8332375, 24'd8020528, 24'd7781523, 24'd7662659, 24'd7687459, 24'd7851015, 24'd8120959, 24'd8443871, 24'd8755846, 
24'd8995145, 24'd9114412, 24'd9090043, 24'd8926862, 24'd8657161, 24'd8334313, 24'd8022211, 24'd7782618, 24'd7662949, 24'd7686886, 24'd7849693, 24'd8119150, 24'd8441932, 24'd8754162, 24'd8994048, 24'd9114120, 24'd9090613, 24'd8928181, 24'd8658969, 24'd8336252, 24'd8023896, 24'd7783716, 24'd7663243, 24'd7686319, 24'd7848375, 24'd8117343, 24'd8439994, 24'd8752475, 24'd8992948, 24'd9113822, 
24'd9091178, 24'd8929497, 24'd8660774, 24'd8338191, 24'd8025584, 24'd7784819, 24'd7663543, 24'd7685756, 24'd7847062, 24'd8115538, 24'd8438055, 24'd8750786, 24'd8991842, 24'd9113520, 24'd9091739, 24'd8930809, 24'd8662579, 24'd8340130, 24'd8027275, 24'd7785927, 24'd7663848, 24'd7685198, 24'd7845752, 24'd8113735, 24'd8436115, 24'd8749094, 24'd8990733, 24'd9113212, 24'd9092294, 24'd8932117, 
24'd8664381, 24'd8342069, 24'd8028968, 24'd7787038, 24'd7664158, 24'd7684645, 24'd7844445, 24'd8111934, 24'd8434176, 24'd8747400, 24'd8989619, 24'd9112900, 24'd9092844, 24'd8933421, 24'd8666181, 24'd8344009, 24'd8030663, 24'd7788154, 24'd7664473, 24'd7684097, 24'd7843143, 24'd8110135, 24'd8432236, 24'd8745703, 24'd8988502, 24'd9112582, 24'd9093390, 24'd8934722, 24'd8667979, 24'd8345949, 
24'd8032361, 24'd7789274, 24'd7664794, 24'd7683555, 24'd7841844, 24'd8108337, 24'd8430296, 24'd8744004, 24'd8987379, 24'd9112259, 24'd9093930, 24'd8936019, 24'd8669776, 24'd8347890, 24'd8034062, 24'd7790398, 24'd7665119, 24'd7683017, 24'd7840549, 24'd8106542, 24'd8428355, 24'd8742302, 24'd8986253, 24'd9111932, 24'd9094466, 24'd8937311, 24'd8671570, 24'd8349830, 24'd8035765, 24'd7791526, 
24'd7665449, 24'd7682483, 24'd7839259, 24'd8104749, 24'd8426414, 24'd8740598, 24'd8985123, 24'd9111599, 24'd9094996, 24'd8938600, 24'd8673362, 24'd8351771, 24'd8037471, 24'd7792659, 24'd7665785, 24'd7681955, 24'd7837971, 24'd8102957, 24'd8424473, 24'd8738891, 24'd8983988, 24'd9111261, 24'd9095522, 24'd8939886, 24'd8675153, 24'd8353713, 24'd8039179, 24'd7793796, 24'd7666125, 24'd7681432, 
24'd7836688, 24'd8101168, 24'd8422532, 24'd8737182, 24'd8982849, 24'd9110918, 24'd9096042, 24'd8941167, 24'd8676941, 24'd8355654, 24'd8040889, 24'd7794937, 24'd7666471, 24'd7680914, 24'd7835409, 24'd8099381, 24'd8420590, 24'd8735470, 24'd8981706, 24'd9110570, 24'd9096558, 24'd8942444, 24'd8678727, 24'd8357596, 24'd8042602, 24'd7796082, 24'd7666821, 24'd7680401, 24'd7834133, 24'd8097595, 
24'd8418648, 24'd8733756, 24'd8980559, 24'd9110217, 24'd9097069, 24'd8943718, 24'd8680512, 24'd8359538, 24'd8044317, 24'd7797231, 24'd7667177, 24'd7679893, 24'd7832862, 24'd8095812, 24'd8416706, 24'd8732039, 24'd8979408, 24'd9109859, 24'd9097575, 24'd8944988, 24'd8682294, 24'd8361480, 24'd8046035, 24'd7798384, 24'd7667537, 24'd7679389, 24'd7831594, 24'd8094031, 24'd8414764, 24'd8730320, 
24'd8978253, 24'd9109495, 24'd9098075, 24'd8946253, 24'd8684074, 24'd8363422, 24'd8047755, 24'd7799542, 24'd7667903, 24'd7678891, 24'd7830330, 24'd8092252, 24'd8412821, 24'd8728599, 24'd8977093, 24'd9109127, 24'd9098571, 24'd8947515, 24'd8685852, 24'd8365365, 24'd8049477, 24'd7800703, 24'd7668274, 24'd7678398, 24'd7829070, 24'd8090475, 24'd8410879, 24'd8726875, 24'd8975929, 24'd9108754, 
24'd9099062, 24'd8948773, 24'd8687628, 24'd8367308, 24'd8051202, 24'd7801869, 24'd7668650, 24'd7677909, 24'd7827815, 24'd8088700, 24'd8408936, 24'd8725149, 24'd8974762, 24'd9108375, 24'd9099548, 24'd8950027, 24'd8689402, 24'd8369250, 24'd8052930, 24'd7803039, 24'd7669031, 24'd7677426, 24'd7826563, 24'd8086927, 24'd8406993, 24'd8723421, 24'd8973590, 24'd9107992, 24'd9100029, 24'd8951277, 
24'd8691174, 24'd8371193, 24'd8054659, 24'd7804213, 24'd7669417, 24'd7676948, 24'd7825314, 24'd8085156, 24'd8405050, 24'd8721690, 24'd8972414, 24'd9107603, 24'd9100505, 24'd8952523, 24'd8692944, 24'd8373136, 24'd8056391, 24'd7805391, 24'd7669808, 24'd7676474, 24'd7824070, 24'd8083387, 24'd8403107, 24'd8719957, 24'd8971234, 24'd9107210, 24'd9100976, 24'd8953765, 24'd8694711, 24'd8375080, 
24'd8058125, 24'd7806573, 24'd7670204, 24'd7676006, 24'd7822830, 24'd8081621, 24'd8401164, 24'd8718222, 24'd8970050, 24'd9106811, 24'd9101442, 24'd8955003, 24'd8696477, 24'd8377023, 24'd8059862, 24'd7807759, 24'd7670605, 24'd7675542, 24'd7821594, 24'd8079857, 24'd8399220, 24'd8716484, 24'd8968861, 24'd9106408, 24'd9101903, 24'd8956238, 24'd8698240, 24'd8378966, 24'd8061601, 24'd7808949, 
24'd7671011, 24'd7675084, 24'd7820362, 24'd8078094, 24'd8397277, 24'd8714744, 24'd8967669, 24'd9105999, 24'd9102358, 24'd8957468, 24'd8700001, 24'd8380910, 24'd8063342, 24'd7810144, 24'd7671422, 24'd7674631, 24'd7819133, 24'd8076334, 24'd8395333, 24'd8713002, 24'd8966473, 24'd9105585, 24'd9102809, 24'd8958694, 24'd8701760, 24'd8382853, 24'd8065085, 24'd7811342, 24'd7671838, 24'd7674182, 
24'd7817909, 24'd8074577, 24'd8393390, 24'd8711257, 24'd8965272, 24'd9105167, 24'd9103255, 24'd8959916, 24'd8703517, 24'd8384797, 24'd8066831, 24'd7812545, 24'd7672260, 24'd7673739, 24'd7816689, 24'd8072821, 24'd8391446, 24'd8709510, 24'd8964068, 24'd9104743, 24'd9103696, 24'd8961135, 24'd8705271, 24'd8386740, 24'd8068579, 24'd7813751, 24'd7672686, 24'd7673300, 24'd7815473, 24'd8071067, 
24'd8389503, 24'd8707761, 24'd8962859, 24'd9104314, 24'd9104132, 24'd8962349, 24'd8707023, 24'd8388684, 24'd8070329, 24'd7814962, 24'd7673117, 24'd7672867, 24'd7814261, 24'd8069316, 24'd8387559, 24'd8706010, 24'd8961647, 24'd9103880, 24'd9104563, 24'd8963559, 24'd8708773, 24'd8390628, 24'd8072082, 24'd7816176, 24'd7673553, 24'd7672439, 24'd7813052, 24'd8067567, 24'd8385616, 24'd8704256, 
24'd8960430, 24'd9103442, 24'd9104989, 24'd8964765, 24'd8710521, 24'd8392571, 24'd8073837, 24'd7817395, 24'd7673995, 24'd7672015, 24'd7811848, 24'd8065821, 24'd8383672, 24'd8702500, 24'd8959210, 24'd9102998, 24'd9105409, 24'd8965967, 24'd8712267, 24'd8394515, 24'd8075593, 24'd7818617, 24'd7674441, 24'd7671597, 24'd7810648, 24'd8064076, 24'd8381729, 24'd8700742, 24'd8957985, 24'd9102549, 
24'd9105825, 24'd8967165, 24'd8714010, 24'd8396458, 24'd8077353, 24'd7819844, 24'd7674892, 24'd7671184, 24'd7809452, 24'd8062334, 24'd8379785, 24'd8698982, 24'd8956756, 24'd9102095, 24'd9106236, 24'd8968359, 24'd8715751, 24'd8398402, 24'd8079114, 24'd7821074, 24'd7675349, 24'd7670775, 24'd7808260, 24'd8060594, 24'd8377842, 24'd8697220, 24'd8955524, 24'd9101636, 24'd9106642, 24'd8969549, 
24'd8717490, 24'd8400345, 24'd8080877, 24'd7822309, 24'd7675810, 24'd7670372, 24'd7807072, 24'd8058857, 24'd8375898, 24'd8695455, 24'd8954287, 24'd9101173, 24'd9107042, 24'd8970735, 24'd8719226, 24'd8402288, 24'd8082643, 24'd7823547, 24'd7676276, 24'd7669974, 24'd7805888, 24'd8057121, 24'd8373955, 24'd8693689, 24'd8953047, 24'd9100704, 24'd9107438, 24'd8971917, 24'd8720960, 24'd8404231, 
24'd8084411, 24'd7824790, 24'd7676747, 24'd7669581, 24'd7804708, 24'd8055389, 24'd8372012, 24'd8691920, 24'd8951802, 24'd9100230, 24'd9107829, 24'd8973095, 24'd8722692, 24'd8406174, 24'd8086180, 24'd7826036, 24'd7677224, 24'd7669193, 24'd7803533, 24'd8053658, 24'd8370069, 24'd8690149, 24'd8950554, 24'd9099751, 24'd9108214, 24'd8974268, 24'd8724421, 24'd8408117, 24'd8087952, 24'd7827287, 
24'd7677705, 24'd7668810, 24'd7802361, 24'd8051930, 24'd8368126, 24'd8688376, 24'd8949302, 24'd9099267, 24'd9108595, 24'd8975438, 24'd8726149, 24'd8410060, 24'd8089727, 24'd7828541, 24'd7678191, 24'd7668432, 24'd7801194, 24'd8050204, 24'd8366183, 24'd8686601, 24'd8948046, 24'd9098779, 24'd9108970, 24'd8976603, 24'd8727873, 24'd8412003, 24'd8091503, 24'd7829799, 24'd7678683, 24'd7668059, 
24'd7800030, 24'd8048480, 24'd8364241, 24'd8684823, 24'd8946785, 24'd9098285, 24'd9109341, 24'd8977765, 24'd8729596, 24'd8413945, 24'd8093281, 24'd7831061, 24'd7679179, 24'd7667691, 24'd7798871, 24'd8046759, 24'd8362298, 24'd8683044, 24'd8945521, 24'd9097786, 24'd9109706, 24'd8978922, 24'd8731315, 24'd8415888, 24'd8095061, 24'd7832327, 24'd7679680, 24'd7667328, 24'd7797716, 24'd8045041, 
24'd8360356, 24'd8681263, 24'd8944253, 24'd9097283, 24'd9110066, 24'd8980075, 24'd8733033, 24'd8417830, 24'd8096844, 24'd7833597, 24'd7680186, 24'd7666970, 24'd7796565, 24'd8043324, 24'd8358414, 24'd8679479, 24'd8942981, 24'd9096774, 24'd9110422, 24'd8981224, 24'd8734748, 24'd8419772, 24'd8098628, 24'd7834871, 24'd7680697, 24'd7666618, 24'd7795418, 24'd8041610, 24'd8356472, 24'd8677694, 
24'd8941706, 24'd9096260, 24'd9110772, 24'd8982368, 24'd8736461, 24'd8421714, 24'd8100415, 24'd7836149, 24'd7681213, 24'd7666270, 24'd7794276, 24'd8039899, 24'd8354531, 24'd8675906, 24'd8940426, 24'd9095742, 24'd9111117, 24'd8983509, 24'd8738171, 24'd8423655, 24'd8102203, 24'd7837430, 24'd7681734, 24'd7665927, 24'd7793137, 24'd8038190, 24'd8352589, 24'd8674117, 24'd8939142, 24'd9095218, 
24'd9111457, 24'd8984645, 24'd8739879, 24'd8425596, 24'd8103994, 24'd7838716, 24'd7682260, 24'd7665590, 24'd7792003, 24'd8036483, 24'd8350648, 24'd8672325, 24'd8937855, 24'd9094690, 24'd9111792, 24'd8985778, 24'd8741584, 24'd8427537, 24'd8105786, 24'd7840005, 24'd7682791, 24'd7665257, 24'd7790873, 24'd8034779, 24'd8348707, 24'd8670532, 24'd8936564, 24'd9094156, 24'd9112122, 24'd8986906, 
24'd8743287, 24'd8429478, 24'd8107581, 24'd7841298, 24'd7683327, 24'd7664930, 24'd7789747, 24'd8033078, 24'd8346767, 24'd8668736, 24'd8935269, 24'd9093618, 24'd9112447, 24'd8988029, 24'd8744987, 24'd8431418, 24'd8109377, 24'd7842595, 24'd7683868, 24'd7664608, 24'd7788625, 24'd8031378, 24'd8344827, 24'd8666939, 24'd8933970, 24'd9093075, 24'd9112767, 24'd8989149, 24'd8746685, 24'd8433358, 
24'd8111176, 24'd7843896, 24'd7684414, 24'd7664290, 24'd7787508, 24'd8029682, 24'd8342887, 24'd8665139, 24'd8932667, 24'd9092526, 24'd9113081, 24'd8990264, 24'd8748381, 24'd8435298, 24'd8112976, 24'd7845201, 24'd7684965, 24'd7663978, 24'd7786395, 24'd8027988, 24'd8340947, 24'd8663338, 24'd8931360, 24'd9091973, 24'd9113391, 24'd8991376, 24'd8750073, 24'd8437238, 24'd8114778, 24'd7846509, 
24'd7685520, 24'd7663671, 24'd7785285, 24'd8026296, 24'd8339008, 24'd8661535, 24'd8930050, 24'd9091415, 24'd9113696, 24'd8992482, 24'd8751764, 24'd8439177, 24'd8116583, 24'd7847821, 24'd7686081, 24'd7663369, 24'd7784181, 24'd8024607, 24'd8337069, 24'd8659730, 24'd8928736, 24'd9090852, 24'd9113995, 24'd8993585, 24'd8753451, 24'd8441116, 24'd8118389, 24'd7849138, 24'd7686646, 24'd7663072, 
24'd7783080, 24'd8022921, 24'd8335130, 24'd8657923, 24'd8927418, 24'd9090284, 24'd9114289, 24'd8994684, 24'd8755137, 24'd8443054, 24'd8120197, 24'd7850457, 24'd7687217, 24'd7662780, 24'd7781984, 24'd8021237, 24'd8333192, 24'd8656114, 24'd8926096, 24'd9089711, 24'd9114579, 24'd8995778, 24'd8756819, 24'd8444992, 24'd8122007, 24'd7851781, 24'd7687792, 24'd7662494, 24'd7780892, 24'd8019555, 
24'd8331254, 24'd8654303, 24'd8924771, 24'd9089133, 24'd9114863, 24'd8996868, 24'd8758499, 24'd8446930, 24'd8123818, 24'd7853108, 24'd7688373, 24'd7662212, 24'd7779804, 24'd8017877, 24'd8329317, 24'd8652490, 24'd8923442, 24'd9088550, 24'd9115142, 24'd8997954, 24'd8760177, 24'd8448867, 24'd8125632, 24'd7854439, 24'd7688958, 24'd7661935, 24'd7778720, 24'd8016201, 24'd8327380, 24'd8650675, 
24'd8922109, 24'd9087963, 24'd9115416, 24'd8999035, 24'd8761852, 24'd8450804, 24'd8127448, 24'd7855774, 24'd7689548, 24'd7661664, 24'd7777641, 24'd8014527, 24'd8325443, 24'd8648859, 24'd8920772, 24'd9087370, 24'd9115685, 24'd9000112, 24'd8763524, 24'd8452740, 24'd8129265, 24'd7857113, 24'd7690143, 24'd7661398, 24'd7776566, 24'd8012856, 24'd8323507, 24'd8647041, 24'd8919431, 24'd9086773, 
24'd9115949, 24'd9001185, 24'd8765193, 24'd8454676, 24'd8131084, 24'd7858455, 24'd7690743, 24'd7661136, 24'd7775495, 24'd8011188, 24'd8321571, 24'd8645221, 24'd8918087, 24'd9086171, 24'd9116207, 24'd9002254, 24'd8766860, 24'd8456612, 24'd8132905, 24'd7859801, 24'd7691347, 24'd7660880, 24'd7774429, 24'd8009522, 24'd8319636, 24'd8643399, 24'd8916739, 24'd9085563, 24'd9116461, 24'd9003318, 
24'd8768525, 24'd8458547, 24'd8134728, 24'd7861151, 24'd7691957, 24'd7660629, 24'd7773367, 24'd8007859, 24'd8317701, 24'd8641575, 24'd8915388, 24'd9084951, 24'd9116710, 24'd9004378, 24'd8770186, 24'd8460481, 24'd8136552, 24'd7862504, 24'd7692572, 24'd7660383, 24'd7772309, 24'd8006199, 24'd8315767, 24'd8639750, 24'd8914032, 24'd9084334, 24'd9116953, 24'd9005433, 24'd8771845, 24'd8462415, 
24'd8138378, 24'd7863862, 24'd7693191, 24'd7660142, 24'd7771255, 24'd8004541, 24'd8313833, 24'd8637923, 24'd8912673, 24'd9083712, 24'd9117191, 24'd9006485, 24'd8773502, 24'd8464348, 24'd8140206, 24'd7865222, 24'd7693815, 24'd7659907, 24'd7770206, 24'd8002886, 24'd8311900, 24'd8636094, 24'd8911311, 24'd9083086, 24'd9117424, 24'd9007532, 24'd8775155, 24'd8466281, 24'd8142036, 24'd7866587, 
24'd7694445, 24'd7659676, 24'd7769161, 24'd8001234, 24'd8309967, 24'd8634263, 24'd8909944, 24'd9082454, 24'd9117652, 24'd9008574, 24'd8776806, 24'd8468214, 24'd8143868, 24'd7867955, 24'd7695079, 24'd7659450, 24'd7768121, 24'd7999585, 24'd8308035, 24'd8632431, 24'd8908574, 24'd9081817, 24'd9117875, 24'd9009613, 24'd8778454, 24'd8470146, 24'd8145701, 24'd7869327, 24'd7695718, 24'd7659230, 
24'd7767085, 24'd7997938, 24'd8306104, 24'd8630597, 24'd8907201, 24'd9081176, 24'd9118093, 24'd9010647, 24'd8780100, 24'd8472077, 24'd8147536, 24'd7870702, 24'd7696361, 24'd7659015, 24'd7766053, 24'd7996294, 24'd8304173, 24'd8628761, 24'd8905824, 24'd9080530, 24'd9118306, 24'd9011676, 24'd8781742, 24'd8474008, 24'd8149372, 24'd7872081, 24'd7697010, 24'd7658804, 24'd7765026, 24'd7994653, 
24'd8302242, 24'd8626924, 24'd8904443, 24'd9079879, 24'd9118514, 24'd9012701, 24'd8783382, 24'd8475938, 24'd8151211, 24'd7873464, 24'd7697663, 24'd7658599, 24'd7764003, 24'd7993014, 24'd8300313, 24'd8625085, 24'd8903058, 24'd9079223, 24'd9118716, 24'd9013722, 24'd8785019, 24'd8477867, 24'd8153051, 24'd7874850, 24'd7698322, 24'd7658399, 24'd7762984, 24'd7991378, 24'd8298383, 24'd8623244, 
24'd8901670, 24'd9078562, 24'd9118914, 24'd9014739, 24'd8786654, 24'd8479796, 24'd8154892, 24'd7876240, 24'd7698985, 24'd7658205, 24'd7761970, 24'd7989745, 24'd8296455, 24'd8621401, 24'd8900278, 24'd9077897, 24'd9119106, 24'd9015751, 24'd8788285, 24'd8481724, 24'd8156735, 24'd7877634, 24'd7699653, 24'd7658015, 24'd7760960, 24'd7988115, 24'd8294527, 24'd8619557, 24'd8898883, 24'd9077226, 
24'd9119293, 24'd9016758, 24'd8789914, 24'd8483652, 24'd8158580, 24'd7879031, 24'd7700326, 24'd7657830, 24'd7759954, 24'd7986488, 24'd8292600, 24'd8617712, 24'd8897484, 24'd9076551, 24'd9119475, 24'd9017762, 24'd8791540, 24'd8485579, 24'd8160427, 24'd7880432, 24'd7701003, 24'd7657651, 24'd7758953, 24'd7984863, 24'd8290673, 24'd8615864, 24'd8896082, 24'd9075871, 24'd9119652, 24'd9018761, 
24'd8793163, 24'd8487505, 24'd8162275, 24'd7881836, 24'd7701686, 24'd7657477, 24'd7757957, 24'd7983241, 24'd8288747, 24'd8614016, 24'd8894676, 24'd9075186, 24'd9119824, 24'd9019755, 24'd8794783, 24'd8489430, 24'd8164125, 24'd7883244, 24'd7702373, 24'd7657307, 24'd7756964, 24'd7981623, 24'd8286822, 24'd8612165, 24'd8893266, 24'd9074496, 24'd9119990, 24'd9020745, 24'd8796401, 24'd8491355, 
24'd8165976, 24'd7884655, 24'd7703065, 24'd7657143, 24'd7755977, 24'd7980007, 24'd8284898, 24'd8610313, 24'd8891853, 24'd9073802, 24'd9120152, 24'd9021731, 24'd8798015, 24'd8493279, 24'd8167829, 24'd7886070, 24'd7703762, 24'd7656984, 24'd7754993, 24'd7978393, 24'd8282974, 24'd8608459, 24'd8890437, 24'd9073103, 24'd9120308, 24'd9022712, 24'd8799627, 24'd8495202, 24'd8169683, 24'd7887488, 
24'd7704464, 24'd7656830, 24'd7754014, 24'd7976783, 24'd8281051, 24'd8606604, 24'd8889016, 24'd9072398, 24'd9120460, 24'd9023688, 24'd8801236, 24'd8497125, 24'd8171539, 24'd7888910, 24'd7705170, 24'd7656682, 24'd7753040, 24'd7975176, 24'd8279129, 24'd8604748, 24'd8887593, 24'd9071690, 24'd9120606, 24'd9024661, 24'd8802842, 24'd8499047, 24'd8173396, 24'd7890335, 24'd7705882, 24'd7656538, 
24'd7752070, 24'd7973571, 24'd8277207, 24'd8602890, 24'd8886166, 24'd9070976, 24'd9120747, 24'd9025628, 24'd8804445, 24'd8500968, 24'd8175255, 24'd7891764, 24'd7706598, 24'd7656400, 24'd7751104, 24'd7971970, 24'd8275287, 24'd8601030, 24'd8884735, 24'd9070257, 24'd9120882, 24'd9026592, 24'd8806045, 24'd8502888, 24'd8177115, 24'd7893197, 24'd7707319, 24'd7656267, 24'd7750143, 24'd7970371, 
24'd8273367, 24'd8599169, 24'd8883301, 24'd9069534, 24'd9121013, 24'd9027551, 24'd8807642, 24'd8504808, 24'd8178977, 24'd7894632, 24'd7708044, 24'd7656138, 24'd7749187, 24'd7968775, 24'd8271448, 24'd8597306, 24'd8881863, 24'd9068806, 24'd9121139, 24'd9028505, 24'd8809236, 24'd8506726, 24'd8180841, 24'd7896072, 24'd7708775, 24'd7656015, 24'd7748235, 24'd7967182, 24'd8269530, 24'd8595442, 
24'd8880422, 24'd9068073, 24'd9121259, 24'd9029455, 24'd8810828, 24'd8508644, 24'd8182706, 24'd7897515, 24'd7709510, 24'd7655897, 24'd7747287, 24'd7965593, 24'd8267612, 24'd8593576, 24'd8878978, 24'd9067336, 24'd9121375, 24'd9030400, 24'd8812416, 24'd8510561, 24'd8184572, 24'd7898961, 24'd7710250, 24'd7655785, 24'd7746344, 24'd7964006, 24'd8265696, 24'd8591710, 24'd8877530, 24'd9066593, 
24'd9121485, 24'd9031341, 24'd8814002, 24'd8512477, 24'd8186440, 24'd7900410, 24'd7710995, 24'd7655677, 24'd7745405, 24'd7962422, 24'd8263780, 24'd8589841, 24'd8876079, 24'd9065846, 24'd9121590, 24'd9032277, 24'd8815584, 24'd8514393, 24'd8188309, 24'd7901863, 24'd7711744, 24'd7655575, 24'd7744471, 24'd7960841, 24'd8261865, 24'd8587971, 24'd8874624, 24'd9065095, 24'd9121690, 24'd9033209, 
24'd8817163, 24'd8516307, 24'd8190179, 24'd7903320, 24'd7712498, 24'd7655477, 24'd7743541, 24'd7959263, 24'd8259951, 24'd8586100, 24'd8873166, 24'd9064338, 24'd9121784, 24'd9034137, 24'd8818740, 24'd8518220, 24'd8192051, 24'd7904780, 24'd7713257, 24'd7655385, 24'd7742616, 24'd7957688, 24'd8258038, 24'd8584228, 24'd8871704, 24'd9063577, 24'd9121874, 24'd9035059, 24'd8820313, 24'd8520133, 
24'd8193924, 24'd7906243, 24'd7714021, 24'd7655298, 24'd7741696, 24'd7956116, 24'd8256126, 24'd8582354, 24'd8870239, 24'd9062811, 24'd9121959, 24'd9035978, 24'd8821883, 24'd8522045, 24'd8195799, 24'd7907710, 24'd7714789, 24'd7655216, 24'd7740780, 24'd7954548, 24'd8254215, 24'd8580478, 24'd8868771, 24'd9062040, 24'd9122038, 24'd9036891, 24'd8823451, 24'd8523955, 24'd8197675, 24'd7909180, 
24'd7715562, 24'd7655139, 24'd7739868, 24'd7952982, 24'd8252305, 24'd8578602, 24'd8867299, 24'd9061264, 24'd9122112, 24'd9037801, 24'd8825015, 24'd8525865, 24'd8199552, 24'd7910653, 24'd7716340, 24'd7655068, 24'd7738961, 24'd7951419, 24'd8250395, 24'd8576724, 24'd8865824, 24'd9060484, 24'd9122181, 24'd9038705, 24'd8826576, 24'd8527774, 24'd8201431, 24'd7912130, 24'd7717123, 24'd7655001, 
24'd7738059, 24'd7949859, 24'd8248487, 24'd8574844, 24'd8864346, 24'd9059699, 24'd9122245, 24'd9039605, 24'd8828134, 24'd8529682, 24'd8203311, 24'd7913610, 24'd7717910, 24'd7654940, 24'd7737161, 24'd7948303, 24'd8246580, 24'd8572964, 24'd8862864, 24'd9058910, 24'd9122304, 24'd9040501, 24'd8829689, 24'd8531589, 24'd8205192, 24'd7915093, 24'd7718702, 24'd7654884, 24'd7736268, 24'd7946749, 
24'd8244673, 24'd8571082, 24'd8861379, 24'd9058115, 24'd9122357, 24'd9041392, 24'd8831241, 24'd8533495, 24'd8207075, 24'd7916580, 24'd7719499, 24'd7654833, 24'd7735379, 24'd7945199, 24'd8242768, 24'd8569198, 24'd8859890, 24'd9057316, 24'd9122406, 24'd9042278, 24'd8832790, 24'd8535399, 24'd8208959, 24'd7918070, 24'd7720300, 24'd7654787, 24'd7734495, 24'd7943651, 24'd8240864, 24'd8567314, 
24'd8858399, 24'd9056513, 24'd9122449, 24'd9043160, 24'd8834336, 24'd8537303, 24'd8210844, 24'd7919563, 24'd7721106, 24'd7654746, 24'd7733616, 24'd7942107, 24'd8238960, 24'd8565428, 24'd8856904, 24'd9055704, 24'd9122487, 24'd9044037, 24'd8835879, 24'd8539206, 24'd8212730, 24'd7921060, 24'd7721917, 24'd7654710, 24'd7732741, 24'd7940566, 24'd8237058, 24'd8563541, 24'd8855405, 24'd9054891, 
24'd9122520, 24'd9044910, 24'd8837418, 24'd8541108, 24'd8214618, 24'd7922560, 24'd7722732, 24'd7654680, 24'd7731871, 24'd7939028, 24'd8235157, 24'd8561653, 24'd8853904, 24'd9054073, 24'd9122548, 24'd9045778, 24'd8838954, 24'd8543008, 24'd8216506, 24'd7924063, 24'd7723552, 24'd7654655, 24'd7731005, 24'd7937494, 24'd8233257, 24'd8559764, 24'd8852399, 24'd9053251, 24'd9122571, 24'd9046641, 
24'd8840488, 24'd8544908, 24'd8218396, 24'd7925569, 24'd7724377, 24'd7654634, 24'd7730144, 24'd7935962, 24'd8231358, 24'd8557873, 24'd8850891, 24'd9052424, 24'd9122589, 24'd9047500, 24'd8842018, 24'd8546806, 24'd8220288, 24'd7927079, 24'd7725206, 24'd7654619, 24'd7729287, 24'd7934434, 24'd8229460, 24'd8555981, 24'd8849380, 24'd9051592, 24'd9122601, 24'd9048354, 24'd8843544, 24'd8548704, 
24'd8222180, 24'd7928592, 24'd7726040, 24'd7654609, 24'd7728435, 24'd7932908, 24'd8227563, 24'd8554088, 24'd8847865, 24'd9050756, 24'd9122609, 24'd9049204, 24'd8845068, 24'd8550600, 24'd8224073, 24'd7930108, 24'd7726879, 24'd7654605, 24'd7727588, 24'd7931386, 24'd8225668, 24'd8552194, 24'd8846348, 24'd9049915, 24'd9122611, 24'd9050049, 24'd8846589, 24'd8552495, 24'd8225968, 24'd7931628, 
24'd7727722, 24'd7654605, 24'd7726746, 24'd7929867, 24'd8223773, 24'd8550299, 24'd8844827, 24'd9049069, 24'd9122608, 24'd9050889, 24'd8848106, 24'd8554389, 24'd8227864, 24'd7933150, 24'd7728570, 24'd7654611, 24'd7725908, 24'd7928352, 24'd8221880, 24'd8548403, 24'd8843302, 24'd9048219, 24'd9122600, 24'd9051724, 24'd8849620, 24'd8556282, 24'd8229761, 24'd7934676, 24'd7729423, 24'd7654621, 
24'd7725074, 24'd7926839, 24'd8219987, 24'd8546505, 24'd8841775, 24'd9047364, 24'd9122586, 24'd9052555, 24'd8851131, 24'd8558173, 24'd8231659, 24'd7936205, 24'd7730280, 24'd7654637, 24'd7724246, 24'd7925330, 24'd8218096, 24'd8544606, 24'd8840245, 24'd9046505, 24'd9122568, 24'd9053382, 24'd8852638, 24'd8560064, 24'd8233558, 24'd7937737, 24'd7731142, 24'd7654658, 24'd7723422, 24'd7923824, 
24'd8216207, 24'd8542707, 24'd8838711, 24'd9045640, 24'd9122544, 24'd9054203, 24'd8854142, 24'd8561953, 24'd8235458, 24'd7939272, 24'd7732008, 24'd7654684, 24'd7722602, 24'd7922322, 24'd8214318, 24'd8540806, 24'd8837174, 24'd9044772, 24'd9122516, 24'd9055020, 24'd8855643, 24'd8563841, 24'd8237360, 24'd7940811, 24'd7732879, 24'd7654716, 24'd7721788, 24'd7920822, 24'd8212431, 24'd8538904, 
24'd8835634, 24'd9043898, 24'd9122482, 24'd9055833, 24'd8857141, 24'd8565728, 24'd8239262, 24'd7942352, 24'd7733755, 24'd7654752, 24'd7720978, 24'd7919326, 24'd8210545, 24'd8537001, 24'd8834091, 24'd9043020, 24'd9122443, 24'd9056640, 24'd8858636, 24'd8567613, 24'd8241166, 24'd7943897, 24'd7734635, 24'd7654794, 24'd7720173, 24'd7917833, 24'd8208660, 24'd8535097, 24'd8832545, 24'd9042138, 
24'd9122399, 24'd9057443, 24'd8860127, 24'd8569497, 24'd8243070, 24'd7945445, 24'd7735520, 24'd7654840, 24'd7719372, 24'd7916344, 24'd8206776, 24'd8533192, 24'd8830995, 24'd9041251, 24'd9122349, 24'd9058242, 24'd8861615, 24'd8571380, 24'd8244976, 24'd7946995, 24'd7736409, 24'd7654892, 24'd7718576, 24'd7914858, 24'd8204894, 24'd8531286, 24'd8829443, 24'd9040359, 24'd9122295, 24'd9059035, 
24'd8863099, 24'd8573262, 24'd8246882, 24'd7948549, 24'd7737303, 24'd7654949, 24'd7717785, 24'd7913375, 24'd8203013, 24'd8529379, 24'd8827887, 24'd9039463, 24'd9122235, 24'd9059824, 24'd8864580, 24'd8575142, 24'd8248790, 24'd7950107, 24'd7738202, 24'd7655011, 24'd7716998, 24'd7911895, 24'd8201133, 24'd8527471, 24'd8826329, 24'd9038562, 24'd9122171, 24'd9060608, 24'd8866058, 24'd8577022, 
24'd8250698, 24'd7951667, 24'd7739105, 24'd7655079, 24'd7716216, 24'd7910419, 24'd8199254, 24'd8525562, 24'd8824767, 24'd9037657, 24'd9122101, 24'd9061388, 24'd8867533, 24'd8578899, 24'd8252608, 24'd7953230, 24'd7740013, 24'd7655151, 24'd7715439, 24'd7908946, 24'd8197377, 24'd8523652, 24'd8823202, 24'd9036747, 24'd9122026, 24'd9062162, 24'd8869004, 24'd8580776, 24'd8254518, 24'd7954796, 
24'd7740925, 24'd7655229, 24'd7714667, 24'd7907477, 24'd8195501, 24'd8521741, 24'd8821635, 24'd9035832, 24'd9121946, 24'd9062932, 24'd8870472, 24'd8582651, 24'd8256429, 24'd7956366, 24'd7741842, 24'd7655311, 24'd7713899, 24'd7906011, 24'd8193627, 24'd8519830, 24'd8820064, 24'd9034913, 24'd9121860, 24'd9063698, 24'd8871936, 24'd8584525, 24'd8258342, 24'd7957938, 24'd7742763, 24'd7655399, 
24'd7713136, 24'd7904548, 24'd8191754, 24'd8517917, 24'd8818490, 24'd9033990, 24'd9121770, 24'd9064458, 24'd8873397, 24'd8586397, 24'd8260255, 24'd7959513, 24'd7743689, 24'd7655492, 24'd7712378, 24'd7903089, 24'd8189882, 24'd8516003, 24'd8816913, 24'd9033062, 24'd9121674, 24'd9065214, 24'd8874855, 24'd8588268, 24'd8262169, 24'd7961092, 24'd7744619, 24'd7655591, 24'd7711625, 24'd7901633, 
24'd8188012, 24'd8514089, 24'd8815333, 24'd9032129, 24'd9121573, 24'd9065965, 24'd8876309, 24'd8590138, 24'd8264084, 24'd7962673, 24'd7745554, 24'd7655694, 24'd7710876, 24'd7900180, 24'd8186143, 24'd8512173, 24'd8813750, 24'd9031192, 24'd9121468, 24'd9066711, 24'd8877760, 24'd8592006, 24'd8266000, 24'd7964257, 24'd7746493, 24'd7655802, 24'd7710132, 24'd7898731, 24'd8184276, 24'd8510257, 
24'd8812164, 24'd9030250, 24'd9121357, 24'd9067453, 24'd8879207, 24'd8593873, 24'd8267916, 24'd7965845, 24'd7747437, 24'd7655916, 24'd7709393, 24'd7897285, 24'd8182410, 24'd8508340, 24'd8810576, 24'd9029304, 24'd9121240, 24'd9068190, 24'd8880651, 24'd8595738, 24'd8269834, 24'd7967435, 24'd7748385, 24'd7656035, 24'd7708659, 24'd7895843, 24'd8180545, 24'd8506422, 24'd8808984, 24'd9028354, 
24'd9121119, 24'd9068922, 24'd8882092, 24'd8597602, 24'd8271752, 24'd7969028, 24'd7749338, 24'd7656158, 24'd7707929, 24'd7894404, 24'd8178682, 24'd8504503, 24'd8807389, 24'd9027399, 24'd9120993, 24'd9069649, 24'd8883529, 24'd8599464, 24'd8273671, 24'd7970624, 24'd7750295, 24'd7656287, 24'd7707204, 24'd7892969, 24'd8176820, 24'd8502584, 24'd8805791, 24'd9026439, 24'd9120861, 24'd9070372, 
24'd8884962, 24'd8601325, 24'd8275591, 24'd7972224, 24'd7751257, 24'd7656421, 24'd7706484, 24'd7891537, 24'd8174960, 24'd8500663, 24'd8804191, 24'd9025475, 24'd9120725, 24'd9071089, 24'd8886392, 24'd8603184, 24'd8277512, 24'd7973826, 24'd7752224, 24'd7656561, 24'd7705769, 24'd7890109, 24'd8173101, 24'd8498742, 24'd8802587, 24'd9024507, 24'd9120583, 24'd9071802, 24'd8887819, 24'd8605042, 
24'd8279434, 24'd7975431, 24'd7753194, 24'd7656705, 24'd7705058, 24'd7888684, 24'd8171244, 24'd8496820, 24'd8800981, 24'd9023534, 24'd9120436, 24'd9072510, 24'd8889242, 24'd8606899, 24'd8281356, 24'd7977038, 24'd7754169, 24'd7656855, 24'd7704352, 24'd7887263, 24'd8169389, 24'd8494897, 24'd8799372, 24'd9022556, 24'd9120284, 24'd9073214, 24'd8890662, 24'd8608754, 24'd8283279, 24'd7978649, 
24'd7755149, 24'd7657009, 24'd7703651, 24'd7885845, 24'd8167535, 24'd8492974, 24'd8797759, 24'd9021575, 24'd9120127, 24'd9073912, 24'd8892078, 24'd8610607, 24'd8285203, 24'd7980263, 24'd7756133, 24'd7657169, 24'd7702955, 24'd7884431, 24'd8165682, 24'd8491050, 24'd8796144, 24'd9020588, 24'd9119964, 24'd9074606, 24'd8893490, 24'd8612459, 24'd8287128, 24'd7981879, 24'd7757122, 24'd7657334, 
24'd7702264, 24'd7883020, 24'd8163831, 24'd8489125, 24'd8794526, 24'd9019598, 24'd9119797, 24'd9075295, 24'd8894899, 24'd8614309, 24'd8289053, 24'd7983499, 24'd7758114, 24'd7657504, 24'd7701577, 24'd7881613, 24'd8161982, 24'd8487199, 24'd8792906, 24'd9018602, 24'd9119624, 24'd9075979, 24'd8896305, 24'd8616158, 24'd8290979, 24'd7985121, 24'd7759112, 24'd7657679, 24'd7700896, 24'd7880209, 
24'd8160134, 24'd8485273, 24'd8791282, 24'd9017603, 24'd9119446, 24'd9076658, 24'd8897706, 24'd8618005, 24'd8292906, 24'd7986746, 24'd7760114, 24'd7657859, 24'd7700219, 24'd7878809, 24'd8158288, 24'd8483346, 24'd8789656, 24'd9016599, 24'd9119264, 24'd9077333, 24'd8899105, 24'd8619850, 24'd8294833, 24'd7988374, 24'd7761120, 24'd7658045, 24'd7699547, 24'd7877413, 24'd8156443, 24'd8481418, 
24'd8788027, 24'd9015591, 24'd9119076, 24'd9078003, 24'd8900499, 24'd8621694, 24'd8296761, 24'd7990004, 24'd7762130, 24'd7658235, 24'd7698879, 24'd7876020, 24'd8154600, 24'd8479490, 24'd8786395, 24'd9014578, 24'd9118883, 24'd9078667, 24'd8901891, 24'd8623536, 24'd8298689, 24'd7991638, 24'd7763145, 24'd7658431, 24'd7698217, 24'd7874630, 24'd8152759, 24'd8477561, 24'd8784760, 24'd9013561, 
24'd9118684, 24'd9079327, 24'd8903278, 24'd8625376, 24'd8300619, 24'd7993274, 24'd7764165, 24'd7658632, 24'd7697559, 24'd7873245, 24'd8150919, 24'd8475631, 24'd8783122, 24'd9012539, 24'd9118481, 24'd9079982, 24'd8904662, 24'd8627215, 24'd8302549, 24'd7994913, 24'd7765188, 24'd7658837, 24'd7696907, 24'd7871862, 24'd8149081, 24'd8473701, 24'd8781482, 24'd9011513, 24'd9118273, 24'd9080633, 
24'd8906042, 24'd8629052, 24'd8304479, 24'd7996554, 24'd7766216, 24'd7659048, 24'd7696259, 24'd7870484, 24'd8147245, 24'd8471771, 24'd8779839, 24'd9010483, 24'd9118059, 24'd9081278, 24'd8907419, 24'd8630888, 24'd8306410, 24'd7998199, 24'd7767249, 24'd7659265, 24'd7695616, 24'd7869109, 24'd8145410, 24'd8469839, 24'd8778193, 24'd9009448, 24'd9117840, 24'd9081919, 24'd8908792, 24'd8632722, 
24'd8308342, 24'd7999846, 24'd7768286, 24'd7659486, 24'd7694978, 24'd7867738, 24'd8143577, 24'd8467907, 24'd8776544, 24'd9008409, 24'd9117617, 24'd9082554, 24'd8910161, 24'd8634554, 24'd8310274, 24'd8001496, 24'd7769327, 24'd7659712, 24'd7694345, 24'd7866370, 24'd8141746, 24'd8465975, 24'd8774893, 24'd9007366, 24'd9117388, 24'd9083185, 24'd8911527, 24'd8636384, 24'd8312207, 24'd8003149, 
24'd7770372, 24'd7659944, 24'd7693716, 24'd7865006, 24'd8139916, 24'd8464042, 24'd8773239, 24'd9006318, 24'd9117154, 24'd9083811, 24'd8912889, 24'd8638213, 24'd8314140, 24'd8004804, 24'd7771422, 24'd7660180, 24'd7693093, 24'd7863646, 24'd8138089, 24'd8462108, 24'd8771582, 24'd9005266, 24'd9116915, 24'd9084432, 24'd8914248, 24'd8640040, 24'd8316074, 24'd8006462, 24'd7772476, 24'd7660422, 
24'd7692474, 24'd7862290, 24'd8136263, 24'd8460174, 24'd8769923, 24'd9004210, 24'd9116670, 24'd9085049, 24'd8915602, 24'd8641865, 24'd8318008, 24'd8008123, 24'd7773535, 24'd7660669, 24'd7691860, 24'd7860937, 24'd8134438, 24'd8458240, 24'd8768261, 24'd9003149, 24'd9116421, 24'd9085660, 24'd8916953, 24'd8643688, 24'd8319943, 24'd8009786, 24'd7774598, 24'd7660920, 24'd7691251, 24'd7859587, 
24'd8132616, 24'd8456305, 24'd8766596, 24'd9002084, 24'd9116167, 24'd9086266, 24'd8918301, 24'd8645510, 24'd8321878, 24'd8011452, 24'd7775665, 24'd7661177, 24'd7690647, 24'd7858242, 24'd8130795, 24'd8454369, 24'd8764929, 24'd9001015, 24'd9115907, 24'd9086868, 24'd8919644, 24'd8647329, 24'd8323814, 24'd8013121, 24'd7776736, 24'd7661440, 24'd7690048, 24'd7856900, 24'd8128976, 24'd8452433, 
24'd8763259, 24'd8999942, 24'd9115643, 24'd9087465, 24'd8920984, 24'd8649147, 24'd8325750, 24'd8014792, 24'd7777812, 24'd7661707, 24'd7689454, 24'd7855562, 24'd8127159, 24'd8450497, 24'd8761586, 24'd8998864, 24'd9115373, 24'd9088056, 24'd8922320, 24'd8650963, 24'd8327687, 24'd8016466, 24'd7778892, 24'd7661979, 24'd7688865, 24'd7854228, 24'd8125344, 24'd8448560, 24'd8759911, 24'd8997782, 
24'd9115098, 24'd9088643, 24'd8923653, 24'd8652778, 24'd8329624, 24'd8018143, 24'd7779976, 24'd7662256, 24'd7688280, 24'd7852897, 24'd8123531, 24'd8446622, 24'd8758233, 24'd8996695, 24'd9114818, 24'd9089225, 24'd8924981, 24'd8654590, 24'd8331561, 24'd8019822, 24'd7781065, 24'd7662539, 24'd7687701, 24'd7851571, 24'd8121719, 24'd8444685, 24'd8756552, 24'd8995605, 24'd9114533, 24'd9089802, 
24'd8926306, 24'd8656401, 24'd8333499, 24'd8021504, 24'd7782157, 24'd7662826, 24'd7687126, 24'd7850248, 24'd8119910, 24'd8442747, 24'd8754869, 24'd8994510, 24'd9114243, 24'd9090374, 24'd8927627, 24'd8658209, 24'd8335438, 24'd8023188, 24'd7783254, 24'd7663119, 24'd7686556, 24'd7848928, 24'd8118102, 24'd8440808, 24'd8753184, 24'd8993411, 24'd9113948, 24'd9090942, 24'd8928945, 24'd8660016, 
24'd8337376, 24'd8024875, 24'd7784356, 24'd7663417, 24'd7685992, 24'd7847613, 24'd8116296, 24'd8438869, 24'd8751496, 24'd8992307, 24'd9113648, 24'd9091504, 24'd8930258, 24'd8661821, 24'd8339315, 24'd8026564, 24'd7785461, 24'd7663719, 24'd7685432, 24'd7846301, 24'd8114492, 24'd8436930, 24'd8749805, 24'd8991200, 24'd9113342, 24'd9092061, 24'd8931568, 24'd8663624, 24'd8341255, 24'd8028256, 
24'd7786571, 24'd7664027, 24'd7684877, 24'd7844994, 24'd8112690, 24'd8434991, 24'd8748112, 24'd8990088, 24'd9113032, 24'd9092614, 24'd8932874, 24'd8665425, 24'd8343194, 24'd8029951, 24'd7787685, 24'd7664340, 24'd7684327, 24'd7843689, 24'd8110890, 24'd8433051, 24'd8746416, 24'd8988972, 24'd9112716, 24'd9093161, 24'd8934176, 24'd8667224, 24'd8345134, 24'd8031648, 24'd7788803, 24'd7664658, 
24'd7683782, 24'd7842389, 24'd8109092, 24'd8431111, 24'd8744718, 24'd8987851, 24'd9112396, 24'd9093704, 24'd8935474, 24'd8669021, 24'd8347075, 24'd8033347, 24'd7789925, 24'd7664982, 24'd7683242, 24'd7841093, 24'd8107296, 24'd8429170, 24'd8743017, 24'd8986727, 24'd9112070, 24'd9094241, 24'd8936769, 24'd8670816, 24'd8349015, 24'd8035049, 24'd7791052, 24'd7665310, 24'd7682707, 24'd7839800, 
24'd8105502, 24'd8427229, 24'd8741314, 24'd8985598, 24'd9111739, 24'd9094774, 24'd8938060, 24'd8672610, 24'd8350956, 24'd8036754, 24'd7792183, 24'd7665643, 24'd7682177, 24'd7838512, 24'd8103710, 24'd8425288, 24'd8739608, 24'd8984465, 24'd9111403, 24'd9095302, 24'd8939346, 24'd8674401, 24'd8352897, 24'd8038461, 24'd7793318, 24'd7665981, 24'd7681651, 24'd7837227, 24'd8101919, 24'd8423347, 
24'd8737900, 24'd8983328, 24'd9111063, 24'd9095824, 24'd8940629, 24'd8676190, 24'd8354839, 24'd8040170, 24'd7794457, 24'd7666325, 24'd7681131, 24'd7835946, 24'd8100131, 24'd8421406, 24'd8736189, 24'd8982187, 24'd9110717, 24'd9096342, 24'd8941908, 24'd8677977, 24'd8356780, 24'd8041882, 24'd7795600, 24'd7666673, 24'd7680616, 24'd7834669, 24'd8098345, 24'd8419464, 24'd8734476, 24'd8981042, 
24'd9110366, 24'd9096855, 24'd8943183, 24'd8679762, 24'd8358722, 24'd8043596, 24'd7796748, 24'd7667027, 24'd7680105, 24'd7833395, 24'd8096561, 24'd8417522, 24'd8732761, 24'd8979892, 24'd9110010, 24'd9097363, 24'd8944455, 24'd8681545, 24'd8360664, 24'd8045313, 24'd7797899, 24'd7667385, 24'd7679600, 24'd7832126, 24'd8094779, 24'd8415580, 24'd8731043, 24'd8978739, 24'd9109648, 24'd9097866, 
24'd8945722, 24'd8683326, 24'd8362607, 24'd8047032, 24'd7799055, 24'd7667749, 24'd7679100, 24'd7830861, 24'd8092999, 24'd8413637, 24'd8729322, 24'd8977581, 24'd9109282, 24'd9098364, 24'd8946986, 24'd8685105, 24'd8364549, 24'd8048754, 24'd7800215, 24'd7668118, 24'd7678604, 24'd7829599, 24'd8091221, 24'd8411695, 24'd8727600, 24'd8976419, 24'd9108911, 24'd9098857, 24'd8948245, 24'd8686882, 
24'd8366492, 24'd8050477, 24'd7801379, 24'd7668491, 24'd7678114, 24'd7828342, 24'd8089445, 24'd8409752, 24'd8725875, 24'd8975253, 24'd9108535, 24'd9099345, 24'd8949501, 24'd8688657, 24'd8368434, 24'd8052204, 24'd7802547, 24'd7668870, 24'd7677628, 24'd7827088, 24'd8087671, 24'd8407809, 24'd8724147, 24'd8974083, 24'd9108153, 24'd9099828, 24'd8950752, 24'd8690430, 24'd8370377, 24'd8053932, 
24'd7803719, 24'd7669254, 24'd7677148, 24'd7825838, 24'd8085900, 24'd8405866, 24'd8722417, 24'd8972908, 24'd9107767, 24'd9100305, 24'd8952000, 24'd8692200, 24'd8372320, 24'd8055663, 24'd7804895, 24'd7669643, 24'd7676672, 24'd7824592, 24'd8084130, 24'd8403923, 24'd8720685, 24'd8971730, 24'd9107376, 24'd9100778, 24'd8953244, 24'd8693969, 24'd8374263, 24'd8057397, 24'd7806076, 24'd7670037, 
24'd7676202, 24'd7823351, 24'd8082363, 24'd8401980, 24'd8718951, 24'd8970547, 24'd9106979, 24'd9101246, 24'd8954484, 24'd8695735, 24'd8376207, 24'd8059132, 24'd7807260, 24'd7670436, 24'd7675736, 24'd7822113, 24'd8080597, 24'd8400037, 24'd8717214, 24'd8969361, 24'd9106578, 24'd9101710, 24'd8955720, 24'd8697499, 24'd8378150, 24'd8060870, 24'd7808449, 24'd7670840, 24'd7675276, 24'd7820879, 
24'd8078834, 24'd8398093, 24'd8715475, 24'd8968170, 24'd9106171, 24'd9102168, 24'd8956952, 24'd8699261, 24'd8380093, 24'd8062610, 24'd7809642, 24'd7671249, 24'd7674820, 24'd7819649, 24'd8077073, 24'd8396150, 24'd8713734, 24'd8966976, 24'd9105760, 24'd9102621, 24'd8958180, 24'd8701021, 24'd8382037, 24'd8064353, 24'd7810838, 24'd7671663, 24'd7674370, 24'd7818423, 24'd8075315, 24'd8394206, 
24'd8711990, 24'd8965777, 24'd9105343, 24'd9103069, 24'd8959403, 24'd8702779, 24'd8383980, 24'd8066098, 24'd7812039, 24'd7672082, 24'd7673924, 24'd7817201, 24'd8073558, 24'd8392263, 24'd8710244, 24'd8964574, 24'd9104921, 24'd9103512, 24'd8960623, 24'd8704534, 24'd8385924, 24'd8067845, 24'd7813244, 24'd7672506, 24'd7673484, 24'd7815983, 24'd8071804, 24'd8390319, 24'd8708496, 24'd8963367, 
24'd9104495, 24'd9103949, 24'd8961839, 24'd8706288, 24'd8387868, 24'd8069594, 24'd7814453, 24'd7672935, 24'd7673048, 24'd7814769, 24'd8070052, 24'd8388376, 24'd8706746, 24'd8962156, 24'd9104063, 24'd9104382, 24'd8963051, 24'd8708039, 24'd8389811, 24'd8071346, 24'd7815665, 24'd7673370, 24'd7672618, 24'd7813559, 24'd8068302, 24'd8386432, 24'd8704993, 24'd8960942, 24'd9103626, 24'd9104810, 
24'd8964259, 24'd8709787, 24'd8391755, 24'd8073099, 24'd7816882, 24'd7673809, 24'd7672193, 24'd7812354, 24'd8066554, 24'd8384489, 24'd8703238, 24'd8959723, 24'd9103185, 24'd9105233, 24'd8965463, 24'd8711534, 24'd8393698, 24'd8074855, 24'd7818103, 24'd7674253, 24'd7671772, 24'd7811152, 24'd8064809, 24'd8382545, 24'd8701481, 24'd8958500, 24'd9102738, 24'd9105651, 24'd8966663, 24'd8713278, 
24'd8395642, 24'd8076613, 24'd7819328, 24'd7674702, 24'd7671357, 24'd7809954, 24'd8063066, 24'd8380601, 24'd8699722, 24'd8957273, 24'd9102286, 24'd9106064, 24'd8967858, 24'd8715020, 24'd8397585, 24'd8078374, 24'd7820557, 24'd7675156, 24'd7670946, 24'd7808760, 24'd8061325, 24'd8378658, 24'd8697960, 24'd8956042, 24'd9101830, 24'd9106472, 24'd8969050, 24'd8716760, 24'd8399529, 24'd8080136, 
24'd7821790, 24'd7675616, 24'd7670541, 24'd7807571, 24'd8059586, 24'd8376715, 24'd8696197, 24'd8954807, 24'd9101368, 24'd9106875, 24'd8970238, 24'd8718497, 24'd8401472, 24'd8081901, 24'd7823027, 24'd7676080, 24'd7670141, 24'd7806385, 24'd8057850, 24'd8374771, 24'd8694431, 24'd8953568, 24'd9100901, 24'd9107273, 24'd8971421, 24'd8720232, 24'd8403415, 24'd8083668, 24'd7824267, 24'd7676549, 
24'd7669745, 24'd7805204, 24'd8056116, 24'd8372828, 24'd8692663, 24'd8952326, 24'd9100430, 24'd9107665, 24'd8972601, 24'd8721965, 24'd8405358, 24'd8085437, 24'd7825512, 24'd7677023, 24'd7669355, 24'd7804026, 24'd8054385, 24'd8370885, 24'd8690893, 24'd8951079, 24'd9099953, 24'd9108053, 24'd8973776, 24'd8723695, 24'd8407301, 24'd8087208, 24'd7826761, 24'd7677502, 24'd7668970, 24'd7802853, 
24'd8052655, 24'd8368942, 24'd8689121, 24'd8949828, 24'd9099471, 24'd9108436, 24'd8974947, 24'd8725423, 24'd8409244, 24'd8088981, 24'd7828014, 24'd7677986, 24'd7668590, 24'd7801684, 24'd8050929, 24'd8366999, 24'd8687346, 24'd8948574, 24'd9098985, 24'd9108813, 24'd8976114, 24'd8727149, 24'd8411187, 24'd8090756, 24'd7829270, 24'd7678476, 24'd7668215, 24'd7800519, 24'd8049204, 24'd8365057, 
24'd8685570, 24'd8947315, 24'd9098493, 24'd9109186, 24'd8977277, 24'd8728872, 24'd8413130, 24'd8092534, 24'd7830531, 24'd7678970, 24'd7667845, 24'd7799358, 24'd8047482, 24'd8363114, 24'd8683792, 24'd8946053, 24'd9097996, 24'd9109553, 24'd8978436, 24'd8730593, 24'd8415072, 24'd8094313, 24'd7831795, 24'd7679469, 24'd7667480, 24'd7798201, 24'd8045762, 24'd8361172, 24'd8682011, 24'd8944786, 
24'd9097495, 24'd9109916, 24'd8979591, 24'd8732312, 24'd8417014, 24'd8096095, 24'd7833063, 24'd7679973, 24'd7667120, 24'd7797048, 24'd8044045, 24'd8359230, 24'd8680229, 24'd8943516, 24'd9096988, 24'd9110273, 24'd8980742, 24'd8734028, 24'd8418956, 24'd8097878, 24'd7834335, 24'd7680482, 24'd7666765, 24'd7795900, 24'd8042330, 24'd8357288, 24'd8678444, 24'd8942242, 24'd9096477, 24'd9110625, 
24'd8981888, 24'd8735742, 24'd8420898, 24'd8099664, 24'd7835612, 24'd7680996, 24'd7666415, 24'd7794755, 24'd8040617, 24'd8355346, 24'd8676657, 24'd8940964, 24'd9095960, 24'd9110973, 24'd8983030, 24'd8737453, 24'd8422840, 24'd8101452, 24'd7836892, 24'd7681515, 24'd7666071, 24'd7793615, 24'd8038907, 24'd8353405, 24'd8674869, 24'd8939682, 24'd9095439, 24'd9111315, 24'd8984168, 24'd8739162, 
24'd8424781, 24'd8103241, 24'd7838175, 24'd7682039, 24'd7665731, 24'd7792479, 24'd8037200, 24'd8351464, 24'd8673078, 24'd8938396, 24'd9094912, 24'd9111652, 24'd8985302, 24'd8740868, 24'd8426722, 24'd8105033, 24'd7839463, 24'd7682568, 24'd7665396, 24'd7791347, 24'd8035495, 24'd8349523, 24'd8671285, 24'd8937107, 24'd9094381, 24'd9111984, 24'd8986432, 24'd8742572, 24'd8428663, 24'd8106827, 
24'd7840755, 24'd7683102, 24'd7665067, 24'd7790219, 24'd8033792, 24'd8347582, 24'd8669491, 24'd8935813, 24'd9093845, 24'd9112311, 24'd8987558, 24'd8744273, 24'd8430603, 24'd8108622, 24'd7842050, 24'd7683640, 24'd7664742, 24'd7789096, 24'd8032092, 24'd8345642, 24'd8667694, 24'd8934516, 24'd9093303, 24'd9112633, 24'd8988679, 24'd8745972, 24'd8432544, 24'd8110420, 24'd7843349, 24'd7684184, 
24'd7664423, 24'd7787977, 24'd8030394, 24'd8343701, 24'd8665895, 24'd8933215, 24'd9092757, 24'd9112950, 24'd8989796, 24'd8747669, 24'd8434484, 24'd8112220, 24'd7844652, 24'd7684733, 24'd7664109, 24'd7786862, 24'd8028699, 24'd8341762, 24'd8664095, 24'd8931910, 24'd9092206, 24'd9113262, 24'd8990909, 24'd8749363, 24'd8436423, 24'd8114021, 24'd7845959, 24'd7685286, 24'd7663799, 24'd7785751, 
24'd8027006, 24'd8339822, 24'd8662292, 24'd8930601, 24'd9091650, 24'd9113568, 24'd8992018, 24'd8751054, 24'd8438362, 24'd8115824, 24'd7847270, 24'd7685845, 24'd7663495, 24'd7784644, 24'd8025316, 24'd8337883, 24'd8660488, 24'd8929288, 24'd9091089, 24'd9113870, 24'd8993122, 24'd8752743, 24'd8440301, 24'd8117630, 24'd7848584, 24'd7686408, 24'd7663196, 24'd7783542, 24'd8023629, 24'd8335944, 
24'd8658682, 24'd8927972, 24'd9090523, 24'd9114166, 24'd8994223, 24'd8754429, 24'd8442240, 24'd8119437, 24'd7849902, 24'd7686977, 24'd7662902, 24'd7782444, 24'd8021944, 24'd8334006, 24'd8656874, 24'd8926652, 24'd9089952, 24'd9114458, 24'd8995319, 24'd8756113, 24'd8444178, 24'd8121246, 24'd7851225, 24'd7687550, 24'd7662613, 24'd7781350, 24'd8020261, 24'd8332068, 24'd8655064, 24'd8925328, 
24'd9089377, 24'd9114744, 24'd8996411, 24'd8757794, 24'd8446116, 24'd8123057, 24'd7852550, 24'd7688128, 24'd7662330, 24'd7780260, 24'd8018582, 24'd8330130, 24'd8653252, 24'd8924000, 24'd9088796, 24'd9115025, 24'd8997498, 24'd8759472, 24'd8448053, 24'd8124870, 24'd7853880, 24'd7688711, 24'd7662051, 24'd7779175, 24'd8016904, 24'd8328193, 24'd8651438, 24'd8922669, 24'd9088210, 24'd9115301, 
24'd8998581, 24'd8761148, 24'd8449990, 24'd8126685, 24'd7855213, 24'd7689299, 24'd7661777, 24'd7778094, 24'd8015230, 24'd8326256, 24'd8649622, 24'd8921334, 24'd9087620, 24'd9115573, 24'd8999660, 24'd8762822, 24'd8451927, 24'd8128501, 24'd7856550, 24'd7689892, 24'd7661509, 24'd7777017, 24'd8013558, 24'd8324320, 24'd8647805, 24'd8919995, 24'd9087024, 24'd9115838, 24'd9000735, 24'd8764492, 
24'd8453863, 24'd8130320, 24'd7857891, 24'd7690490, 24'd7661245, 24'd7775944, 24'd8011888, 24'd8322384, 24'd8645986, 24'd8918652, 24'd9086424, 24'd9116099, 24'd9001805, 24'd8766160, 24'd8455799, 24'd8132140, 24'd7859235, 24'd7691093, 24'd7660987, 24'd7774876, 24'd8010222, 24'd8320449, 24'd8644164, 24'd8917306, 24'd9085819, 24'd9116355, 24'd9002871, 24'd8767826, 24'd8457734, 24'd8133962, 
24'd7860584, 24'd7691700, 24'd7660734, 24'd7773812, 24'd8008557, 24'd8318514, 24'd8642342, 24'd8915956, 24'd9085209, 24'd9116606, 24'd9003933, 24'd8769489, 24'd8459668, 24'd8135785, 24'd7861936, 24'd7692313, 24'd7660486, 24'd7772753, 24'd8006896, 24'd8316579, 24'd8640517, 24'd8914602, 24'd9084594, 24'd9116851, 24'd9004991, 24'd8771149, 24'd8461603, 24'd8137611, 24'd7863291, 24'd7692930, 
24'd7660243, 24'd7771697, 24'd8005237, 24'd8314645, 24'd8638691, 24'd8913245, 24'd9083974, 24'd9117092, 24'd9006044, 24'd8772806, 24'd8463536, 24'd8139438, 24'd7864650, 24'd7693553, 24'd7660005, 24'd7770646, 24'd8003581, 24'd8312712, 24'd8636862, 24'd8911884, 24'd9083349, 24'd9117327, 24'd9007092, 24'd8774461, 24'd8465470, 24'd8141267, 24'd7866013, 24'd7694180, 24'd7659772, 24'd7769600, 
24'd8001928, 24'd8310779, 24'd8635032, 24'd8910519, 24'd9082720, 24'd9117557, 24'd9008137, 24'd8776113, 24'd8467402, 24'd8143098, 24'd7867380, 24'd7694812, 24'd7659544, 24'd7768557, 24'd8000277, 24'd8308847, 24'd8633201, 24'd8909150, 24'd9082085, 24'd9117782, 24'd9009177, 24'd8777762, 24'd8469334, 24'd8144931, 24'd7868750, 24'd7695449, 24'd7659322, 24'd7767519, 24'd7998629, 24'd8306915, 
24'd8631368, 24'd8907778, 24'd9081446, 24'd9118002, 24'd9010213, 24'd8779409, 24'd8471266, 24'd8146765, 24'd7870124, 24'd7696090, 24'd7659104, 24'd7766486, 24'd7996984, 24'd8304984, 24'd8629532, 24'd8906403, 24'd9080802, 24'd9118217, 24'd9011244, 24'd8781053, 24'd8473197, 24'd8148601, 24'd7871502, 24'd7696737, 24'd7658892, 24'd7765457, 24'd7995342, 24'd8303053, 24'd8627696, 24'd8905023, 
24'd9080153, 24'd9118427, 24'd9012271, 24'd8782694, 24'd8475127, 24'd8150438, 24'd7872883, 24'd7697388, 24'd7658685, 24'd7764432, 24'd7993702, 24'd8301123, 24'd8625857, 24'd8903640, 24'd9079499, 24'd9118632, 24'd9013294, 24'd8784332, 24'd8477057, 24'd8152278, 24'd7874268, 24'd7698045, 24'd7658483, 24'd7763411, 24'd7992065, 24'd8299194, 24'd8624017, 24'd8902254, 24'd9078840, 24'd9118831, 
24'd9014312, 24'd8785967, 24'd8478986, 24'd8154118, 24'd7875656, 24'd7698706, 24'd7658286, 24'd7762395, 24'd7990431, 24'd8297265, 24'd8622175, 24'd8900863, 24'd9078177, 24'd9119026, 24'd9015326, 24'd8787600, 24'd8480914, 24'd8155961, 24'd7877048, 24'd7699372, 24'd7658094, 24'd7761384, 24'd7988799, 24'd8295337, 24'd8620332, 24'd8899470, 24'd9077508, 24'd9119215, 24'd9016336, 24'd8789230, 
24'd8482842, 24'd8157805, 24'd7878444, 24'd7700043, 24'd7657907, 24'd7760376, 24'd7987171, 24'd8293409, 24'd8618487, 24'd8898072, 24'd9076835, 24'd9119399, 24'd9017341, 24'd8790857, 24'd8484769, 24'd8159651, 24'd7879843, 24'd7700718, 24'd7657726, 24'd7759373, 24'd7985545, 24'd8291482, 24'd8616641, 24'd8896671, 24'd9076157, 24'd9119578, 24'd9018342, 24'd8792482, 24'd8486696, 24'd8161498, 
24'd7881246, 24'd7701399, 24'd7657549, 24'd7758375, 24'd7983922, 24'd8289556, 24'd8614792, 24'd8895267, 24'd9075474, 24'd9119752, 24'd9019338, 24'd8794103, 24'd8488622, 24'd8163347, 24'd7882652, 24'd7702084, 24'd7657378, 24'd7757381, 24'd7982302, 24'd8287631, 24'd8612943, 24'd8893859, 24'd9074787, 24'd9119921, 24'd9020330, 24'd8795722, 24'd8490547, 24'd8165198, 24'd7884062, 24'd7702774, 
24'd7657212, 24'd7756391, 24'd7980685, 24'd8285706, 24'd8611091, 24'd8892447, 24'd9074094, 24'd9120085, 24'd9021317, 24'd8797338, 24'd8492471, 24'd8167050, 24'd7885475, 24'd7703469, 24'd7657050, 24'd7755406, 24'd7979071, 24'd8283782, 24'd8609238, 24'd8891032, 24'd9073397, 24'd9120243, 24'd9022300, 24'd8798950, 24'd8494395, 24'd8168904, 24'd7886892, 24'd7704169, 24'd7656894, 24'd7754425, 
24'd7977459, 24'd8281859, 24'd8607384, 24'd8889613, 24'd9072695, 24'd9120397, 24'd9023279, 24'd8800560, 24'd8496318, 24'd8170759, 24'd7888312, 24'd7704873, 24'd7656744, 24'd7753449, 24'd7975851, 24'd8279936, 24'd8605528, 24'd8888191, 24'd9071988, 24'd9120545, 24'd9024253, 24'd8802168, 24'd8498240, 24'd8172616, 24'd7889736, 24'd7705582, 24'd7656598, 24'd7752477, 24'd7974245, 24'd8278014, 
24'd8603670, 24'd8886766, 24'd9071276, 24'd9120688, 24'd9025222, 24'd8803772, 24'd8500161, 24'd8174474, 24'd7891164, 24'd7706296, 24'd7656457, 24'd7751509, 24'd7972642, 24'd8276093, 24'd8601811, 24'd8885336, 24'd9070560, 24'd9120826, 24'd9026188, 24'd8805373, 24'd8502082, 24'd8176334, 24'd7892595, 24'd7707015, 24'd7656322, 24'd7750546, 24'd7971042, 24'd8274173, 24'd8599951, 24'd8883904, 
24'd9069839, 24'd9120959, 24'd9027148, 24'd8806972, 24'd8504002, 24'd8178195, 24'd7894029, 24'd7707739, 24'd7656192, 24'd7749588, 24'd7969445, 24'd8272254, 24'd8598089, 24'd8882468, 24'd9069112, 24'd9121087, 24'd9028105, 24'd8808567, 24'd8505921, 24'd8180058, 24'd7895467, 24'd7708467, 24'd7656066, 24'd7748634, 24'd7967851, 24'd8270335, 24'd8596225, 24'd8881028, 24'd9068382, 24'd9121209, 
24'd9029056, 24'd8810160, 24'd8507839, 24'd8181922, 24'd7896908, 24'd7709201, 24'd7655946, 24'd7747684, 24'd7966260, 24'd8268418, 24'd8594360, 24'd8879585, 24'd9067646, 24'd9121327, 24'd9030004, 24'd8811749, 24'd8509756, 24'd8183788, 24'd7898353, 24'd7709938, 24'd7655831, 24'd7746739, 24'd7964672, 24'd8266501, 24'd8592494, 24'd8878139, 24'd9066906, 24'd9121439, 24'd9030946, 24'd8813336, 
24'd8511673, 24'd8185655, 24'd7899801, 24'd7710681, 24'd7655722, 24'd7745799, 24'd7963087, 24'd8264585, 24'd8590626, 24'd8876689, 24'd9066161, 24'd9121546, 24'd9031885, 24'd8814920, 24'd8513588, 24'd8187523, 24'd7901253, 24'd7711429, 24'd7655617, 24'd7744863, 24'd7961505, 24'd8262669, 24'd8588757, 24'd8875235, 24'd9065411, 24'd9121648, 24'd9032818, 24'd8816500, 24'd8515503, 24'd8189393, 
24'd7902708, 24'd7712181, 24'd7655518, 24'd7743931, 24'd7959926, 24'd8260755, 24'd8586886, 24'd8873779, 24'd9064656, 24'd9121745, 24'd9033748, 24'd8818078, 24'd8517417, 24'd8191265, 24'd7904166, 24'd7712938, 24'd7655423, 24'd7743004, 24'd7958349, 24'd8258842, 24'd8585014, 24'd8872318, 24'd9063897, 24'd9121837, 24'd9034672, 24'd8819653, 24'd8519330, 24'd8193137, 24'd7905628, 24'd7713699, 
24'd7655334, 24'd7742082, 24'd7956776, 24'd8256929, 24'd8583141, 24'd8870855, 24'd9063133, 24'd9121924, 24'd9035593, 24'd8821224, 24'd8521242, 24'd8195011, 24'd7907093, 24'd7714466, 24'd7655250, 24'd7741164, 24'd7955206, 24'd8255018, 24'd8581266, 24'd8869388, 24'd9062364, 24'd9122005, 24'd9036508, 24'd8822793, 24'd8523153, 24'd8196887, 24'd7908562, 24'd7715237, 24'd7655171, 24'd7740251, 
24'd7953639, 24'd8253107, 24'd8579390, 24'd8867918, 24'd9061591, 24'd9122082, 24'd9037419, 24'd8824358, 24'd8525063, 24'd8198764, 24'd7910034, 24'd7716013, 24'd7655097, 24'd7739342, 24'd7952075, 24'd8251197, 24'd8577513, 24'd8866444, 24'd9060812, 24'd9122153, 24'd9038326, 24'd8825921, 24'd8526972, 24'd8200642, 24'd7911509, 24'd7716793, 24'd7655029, 24'd7738438, 24'd7950514, 24'd8249288, 
24'd8575634, 24'd8864967, 24'd9060030, 24'd9122219, 24'd9039228, 24'd8827480, 24'd8528881, 24'd8202521, 24'd7912988, 24'd7717579, 24'd7654965, 24'd7737538, 24'd7948956, 24'd8247381, 24'd8573754, 24'd8863487, 24'd9059242, 24'd9122280, 24'd9040125, 24'd8829037, 24'd8530788, 24'd8204402, 24'd7914470, 24'd7718369, 24'd7654907, 24'd7736643, 24'd7947401, 24'd8245474, 24'd8571872, 24'd8862003, 
24'd9058450, 24'd9122336, 24'd9041018, 24'd8830590, 24'd8532694, 24'd8206284, 24'd7915955, 24'd7719163, 24'd7654853, 24'd7735752, 24'd7945850, 24'd8243568, 24'd8569990, 24'd8860516, 24'd9057652, 24'd9122386, 24'd9041906, 24'd8832140, 24'd8534599, 24'd8208167, 24'd7917444, 24'd7719963, 24'd7654805, 24'd7734866, 24'd7944301, 24'd8241663, 24'd8568106, 24'd8859026, 24'd9056851, 24'd9122432, 
24'd9042790, 24'd8833687, 24'd8536504, 24'd8210052, 24'd7918936, 24'd7720767, 24'd7654762, 24'd7733985, 24'd7942756, 24'd8239760, 24'd8566221, 24'd8857532, 24'd9056044, 24'd9122472, 24'd9043669, 24'd8835231, 24'd8538407, 24'd8211938, 24'd7920431, 24'd7721576, 24'd7654725, 24'd7733108, 24'd7941213, 24'd8237857, 24'd8564334, 24'd8856035, 24'd9055233, 24'd9122507, 24'd9044544, 24'd8836772, 
24'd8540309, 24'd8213825, 24'd7921929, 24'd7722389, 24'd7654692, 24'd7732236, 24'd7939674, 24'd8235955, 24'd8562446, 24'd8854535, 24'd9054417, 24'd9122537, 24'd9045414, 24'd8838309, 24'd8542210, 24'd8215713, 24'd7923431, 24'd7723207, 24'd7654665, 24'd7731368, 24'd7938138, 24'd8234055, 24'd8560558, 24'd8853032, 24'd9053597, 24'd9122562, 24'd9046279, 24'd8839844, 24'd8544110, 24'd8217602, 
24'd7924936, 24'd7724030, 24'd7654642, 24'd7730505, 24'd7936605, 24'd8232155, 24'd8558667, 24'd8851525, 24'd9052772, 24'd9122582, 24'd9047140, 24'd8841375, 24'd8546009, 24'd8219493, 24'd7926445, 24'd7724857, 24'd7654625, 24'd7729647, 24'd7935075, 24'd8230257, 24'd8556776, 24'd8850015, 24'd9051942, 24'd9122597, 24'd9047996, 24'd8842904, 24'd8547907, 24'd8221385, 24'd7927956, 24'd7725689, 
24'd7654613, 24'd7728793, 24'd7933549, 24'd8228360, 24'd8554884, 24'd8848502, 24'd9051108, 24'd9122606, 24'd9048847, 24'd8844428, 24'd8549803, 24'd8223278, 24'd7929471, 24'd7726526, 24'd7654606, 24'd7727944, 24'd7932025, 24'd8226464, 24'd8552990, 24'd8846985, 24'd9050269, 24'd9122610, 24'd9049694, 24'd8845950, 24'd8551699, 24'd8225172, 24'd7930989, 24'd7727368, 24'd7654604, 24'd7727099, 
24'd7930505, 24'd8224569, 24'd8551095, 24'd8845466, 24'd9049425, 24'd9122610, 24'd9050536, 24'd8847469, 24'd8553593, 24'd8227068, 24'd7932510, 24'd7728214, 24'd7654608, 24'd7726259, 24'd7928988, 24'd8222675, 24'd8549199, 24'd8843943, 24'd9048577, 24'd9122604, 24'd9051374, 24'd8848984, 24'd8555487, 24'd8228964, 24'd7934035, 24'd7729064, 24'd7654616, 24'd7725424, 24'd7927474, 24'd8220782, 
24'd8547302, 24'd8842417, 24'd9047724, 24'd9122593, 24'd9052207, 24'd8850496, 24'd8557379, 24'd8230862, 24'd7935562, 24'd7729919, 24'd7654630, 24'd7724593, 24'd7925964, 24'd8218891, 24'd8545404, 24'd8840888, 24'd9046866, 24'd9122576, 24'd9053035, 24'd8852005, 24'd8559270, 24'd8232760, 24'd7937093, 24'd7730779, 24'd7654649, 24'd7723767, 24'd7924457, 24'd8217000, 24'd8543505, 24'd8839356, 
24'd9046004, 24'd9122555, 24'd9053859, 24'd8853511, 24'd8561159, 24'd8234660, 24'd7938627, 24'd7731644, 24'd7654673, 24'd7722946, 24'd7922953, 24'd8215111, 24'd8541605, 24'd8837820, 24'd9045137, 24'd9122528, 24'd9054678, 24'd8855013, 24'd8563048, 24'd8236561, 24'd7940164, 24'd7732513, 24'd7654702, 24'd7722129, 24'd7921452, 24'd8213223, 24'd8539703, 24'd8836281, 24'd9044266, 24'd9122497, 
24'd9055492, 24'd8856512, 24'd8564935, 24'd8238463, 24'd7941704, 24'd7733387, 24'd7654736, 24'd7721317, 24'd7919954, 24'd8211337, 24'd8537801, 24'd8834740, 24'd9043390, 24'd9122460, 24'd9056302, 24'd8858008, 24'd8566821, 24'd8240366, 24'd7943248, 24'd7734265, 24'd7654776, 24'd7720510, 24'd7918460, 24'd8209451, 24'd8535897, 24'd8833195, 24'd9042509, 24'd9122418, 24'd9057107, 24'd8859501, 
24'd8568706, 24'd8242270, 24'd7944794, 24'd7735148, 24'd7654820, 24'd7719708, 24'd7916969, 24'd8207567, 24'd8533993, 24'd8831647, 24'd9041624, 24'd9122371, 24'd9057907, 24'd8860990, 24'd8570590, 24'd8244175, 24'd7946344, 24'd7736035, 24'd7654870, 24'd7718910, 24'd7915482, 24'd8205684, 24'd8532087, 24'd8830095, 24'd9040734, 24'd9122318, 24'd9058702, 24'd8862476, 24'd8572472, 24'd8246081, 
24'd7947896, 24'd7736927, 24'd7654925, 24'd7718117, 24'd7913997, 24'd8203803, 24'd8530180, 24'd8828541, 24'd9039840, 24'd9122261, 24'd9059493, 24'd8863959, 24'd8574353, 24'd8247988, 24'd7949452, 24'd7737824, 24'd7654985, 24'd7717328, 24'd7912516, 24'd8201922, 24'd8528273, 24'd8826984, 24'd9038941, 24'd9122198, 24'd9060279, 24'd8865438, 24'd8576232, 24'd8249896, 24'd7951011, 24'd7738725, 
24'd7655050, 24'd7716544, 24'd7911039, 24'd8200043, 24'd8526364, 24'd8825423, 24'd9038038, 24'd9122131, 24'd9061061, 24'd8866914, 24'd8578111, 24'd8251805, 24'd7952573, 24'd7739631, 24'd7655120, 24'd7715765, 24'd7909565, 24'd8198166, 24'd8524455, 24'd8823860, 24'd9037130, 24'd9122058, 24'd9061838, 24'd8868386, 24'd8579988, 24'd8253715, 24'd7954138, 24'd7740541, 24'd7655196, 24'd7714991, 
24'd7908094, 24'd8196289, 24'd8522544, 24'd8822293, 24'd9036217, 24'd9121980, 24'd9062610, 24'd8869856, 24'd8581863, 24'd8255626, 24'd7955706, 24'd7741456, 24'd7655276, 24'd7714221, 24'd7906626, 24'd8194414, 24'd8520633, 24'd8820724, 24'd9035300, 24'd9121897, 24'd9063377, 24'd8871321, 24'd8583738, 24'd8257538, 24'd7957277, 24'd7742375, 24'd7655362, 24'd7713456, 24'd7905162, 24'd8192541, 
24'd8518721, 24'd8819151, 24'd9034378, 24'd9121808, 24'd9064139, 24'd8872784, 24'd8585611, 24'd8259451, 24'd7958851, 24'd7743299, 24'd7655453, 24'd7712696, 24'd7903701, 24'd8190668, 24'd8516807, 24'd8817576, 24'd9033452, 24'd9121715, 24'd9064897, 24'd8874243, 24'd8587482, 24'd8261365, 24'd7960428, 24'd7744228, 24'd7655549, 24'd7711941, 24'd7902244, 24'd8188797, 24'd8514893, 24'd8815997, 
24'd9032521, 24'd9121616, 24'd9065650, 24'd8875699, 24'd8589352, 24'd8263279, 24'd7962008, 24'd7745161, 24'd7655650, 24'd7711190, 24'd7900790, 24'd8186928, 24'd8512978, 24'd8814415, 24'd9031586, 24'd9121513, 24'd9066399, 24'd8877151, 24'd8591221, 24'd8265195, 24'd7963591, 24'd7746098, 24'd7655756, 24'd7710444, 24'd7899339, 24'd8185060, 24'd8511062, 24'd8812831, 24'd9030647, 24'd9121404, 
24'd9067142, 24'd8878600, 24'd8593089, 24'd8267111, 24'd7965178, 24'd7747040, 24'd7655867, 24'd7709703, 24'd7897892, 24'd8183193, 24'd8509145, 24'd8811243, 24'd9029702, 24'd9121290, 24'd9067881, 24'd8880045, 24'd8594955, 24'd8269028, 24'd7966767, 24'd7747986, 24'd7655984, 24'd7708966, 24'd7896449, 24'd8181328, 24'd8507228, 24'd8809653, 24'd9028754, 24'd9121171, 24'd9068615, 24'd8881487, 
24'd8596819, 24'd8270946, 24'd7968359, 24'd7748937, 24'd7656106, 24'd7708235, 24'd7895008, 24'd8179464, 24'd8505309, 24'd8808059, 24'd9027800, 24'd9121047, 24'd9069344, 24'd8882925, 24'd8598682, 24'd8272865, 24'd7969954, 24'd7749893, 24'd7656233, 24'd7707508, 24'd7893572, 24'd8177602, 24'd8503390, 24'd8806463, 24'd9026843, 24'd9120917, 24'd9070069, 24'd8884360, 24'd8600544, 24'd8274785, 
24'd7971551, 24'd7750853, 24'd7656364, 24'd7706786, 24'd7892138, 24'd8175741, 24'd8501470, 24'd8804863, 24'd9025881, 24'd9120783, 24'd9070788, 24'd8885792, 24'd8602404, 24'd8276705, 24'd7973152, 24'd7751817, 24'd7656502, 24'd7706068, 24'd7890709, 24'd8173882, 24'd8499549, 24'd8803261, 24'd9024914, 24'd9120643, 24'd9071503, 24'd8887220, 24'd8604262, 24'd8278627, 24'd7974756, 24'd7752786, 
24'd7656644, 24'd7705356, 24'd7889282, 24'd8172024, 24'd8497628, 24'd8801656, 24'd9023943, 24'd9120498, 24'd9072214, 24'd8888645, 24'd8606119, 24'd8280549, 24'd7976363, 24'd7753759, 24'd7656791, 24'd7704648, 24'd7887859, 24'd8170168, 24'd8495705, 24'd8800048, 24'd9022967, 24'd9120348, 24'd9072919, 24'd8890066, 24'd8607975, 24'd8282471, 24'd7977972, 24'd7754737, 24'd7656944, 24'd7703945, 
24'd7886440, 24'd8168313, 24'd8493782, 24'd8798437, 24'd9021987, 24'd9120193, 24'd9073620, 24'd8891483, 24'd8609829, 24'd8284395, 24'd7979585, 24'd7755719, 24'd7657101, 24'd7703247, 24'd7885024, 24'd8166460, 24'd8491858, 24'd8796823, 24'd9021003, 24'd9120033, 24'd9074315, 24'd8892897, 24'd8611681, 24'd8286319, 24'd7981200, 24'd7756706, 24'd7657264, 24'd7702554, 24'd7883612, 24'd8164608, 
24'd8489933, 24'd8795206, 24'd9020014, 24'd9119868, 24'd9075006, 24'd8894308, 24'd8613532, 24'd8288244, 24'd7982818, 24'd7757697, 24'd7657432, 24'd7701865, 24'd7882203, 24'd8162758, 24'd8488008, 24'd8793587, 24'd9019021, 24'd9119697, 24'd9075692, 24'd8895715, 24'd8615381, 24'd8290170, 24'd7984439, 24'd7758692, 24'd7657605, 24'd7701181, 24'd7880798, 24'd8160910, 24'd8486082, 24'd8791964, 
24'd9018023, 24'd9119522, 24'd9076374, 24'd8897118, 24'd8617229, 24'd8292096, 24'd7986063, 24'd7759692, 24'd7657783, 24'd7700502, 24'd7879397, 24'd8159063, 24'd8484155, 24'd8790339, 24'd9017021, 24'd9119341, 24'd9077050, 24'd8898518, 24'd8619075, 24'd8294023, 24'd7987689, 24'd7760697, 24'd7657966, 24'd7699828, 24'd7877999, 24'd8157218, 24'd8482228, 24'd8788711, 24'd9016015, 24'd9119155, 
24'd9077722, 24'd8899914, 24'd8620919, 24'd8295951, 24'd7989319, 24'd7761705, 24'd7658155, 24'd7699159, 24'd7876604, 24'd8155374, 24'd8480300, 24'd8787080, 24'd9015004, 24'd9118964, 24'd9078389, 24'd8901307, 24'd8622762, 24'd8297879, 24'd7990951, 24'd7762718, 24'd7658348, 24'd7698495, 24'd7875213, 24'd8153532, 24'd8478371, 24'd8785447, 24'd9013988, 24'd9118768, 24'd9079051, 24'd8902696, 
24'd8624604, 24'd8299808, 24'd7992586, 24'd7763736, 24'd7658547, 24'd7697835, 24'd7873826, 24'd8151691, 24'd8476442, 24'd8783810, 24'd9012969, 24'd9118567, 24'd9079708, 24'd8904081, 24'd8626443, 24'd8301738, 24'd7994224, 24'd7764758, 24'd7658750, 24'd7697180, 24'd7872443, 24'd8149853, 24'd8474512, 24'd8782171, 24'd9011945, 24'd9118361, 24'd9080360, 24'd8905463, 24'd8628281, 24'd8303668, 
24'd7995864, 24'd7765784, 24'd7658959, 24'd7696530, 24'd7871062, 24'd8148016, 24'd8472582, 24'd8780529, 24'd9010916, 24'd9118149, 24'd9081008, 24'd8906841, 24'd8630117, 24'd8305599, 24'd7997508, 24'd7766815, 24'd7659173, 24'd7695885, 24'd7869686, 24'd8146180, 24'd8470650, 24'd8778884, 24'd9009883, 24'd9117933, 24'd9081650, 24'd8908216, 24'd8631952, 24'd8307530, 24'd7999154, 24'd7767850, 
24'd7659392, 24'd7695245, 24'd7868313, 24'd8144347, 24'd8468719, 24'd8777237, 24'd9008846, 24'd9117711, 24'd9082288, 24'd8909587, 24'd8633784, 24'd8309462, 24'd8000803, 24'd7768889, 24'd7659616, 24'd7694610, 24'd7866944, 24'd8142515, 24'd8466787, 24'd8775587, 24'd9007805, 24'd9117485, 24'd9082921, 24'd8910954, 24'd8635616, 24'd8311395, 24'd8002454, 24'd7769933, 24'd7659846, 24'd7693979, 
24'd7865579, 24'd8140685, 24'd8464854, 24'd8773934, 24'd9006759, 24'd9117253, 24'd9083549, 24'd8912318, 24'd8637445, 24'd8313328, 24'd8004108, 24'd7770981, 24'd7660080, 24'd7693354, 24'd7864217, 24'd8138856, 24'd8462920, 24'd8772278, 24'd9005709, 24'd9117016, 24'd9084172, 24'd8913678, 24'd8639273, 24'd8315261, 24'd8005765, 24'd7772033, 24'd7660320, 24'd7692733, 24'd7862859, 24'd8137029, 
24'd8460987, 24'd8770620, 24'd9004654, 24'd9116774, 24'd9084790, 24'd8915034, 24'd8641098, 24'd8317196, 24'd8007425, 24'd7773090, 24'd7660564, 24'd7692117, 24'd7861504, 24'd8135204, 24'd8459052, 24'd8768959, 24'd9003595, 24'd9116526, 24'd9085404, 24'd8916386, 24'd8642922, 24'd8319130, 24'd8009087, 24'd7774151, 24'd7660814, 24'd7691506, 24'd7860154, 24'd8133381, 24'd8457117, 24'd8767296, 
24'd9002532, 24'd9116274, 24'd9086012, 24'd8917735, 24'd8644745, 24'd8321065, 24'd8010752, 24'd7775216, 24'd7661069, 24'd7690900, 24'd7858807, 24'd8131560, 24'd8455182, 24'd8765629, 24'd9001465, 24'd9116017, 24'd9086616, 24'd8919080, 24'd8646565, 24'd8323001, 24'd8012420, 24'd7776286, 24'd7661329, 24'd7690299, 24'd7857463, 24'd8129740, 24'd8453246, 24'd8763960, 24'd9000393, 24'd9115754, 
24'd9087215, 24'd8920422, 24'd8648384, 24'd8324937, 24'd8014090, 24'd7777359, 24'd7661594, 24'd7689703, 24'd7856124, 24'd8127922, 24'd8451310, 24'd8762289, 24'd8999317, 24'd9115487, 24'd9087808, 24'd8921760, 24'd8650201, 24'd8326873, 24'd8015763, 24'd7778438, 24'd7661864, 24'd7689112, 24'd7854788, 24'd8126106, 24'd8449373, 24'd8760615, 24'd8998237, 24'd9115214, 24'd9088397, 24'd8923094, 
24'd8652016, 24'd8328810, 24'd8017438, 24'd7779520, 24'd7662139, 24'd7688525, 24'd7853456, 24'd8124292, 24'd8447436, 24'd8758938, 24'd8997152, 24'd9114936, 24'd9088981, 24'd8924424, 24'd8653829, 24'd8330748, 24'd8019116, 24'd7780607, 24'd7662420, 24'd7687943, 24'd7852128, 24'd8122480, 24'd8445499, 24'd8757259, 24'd8996063, 24'd9114653, 24'd9089560, 24'd8925750, 24'd8655640, 24'd8332685, 
24'd8020797, 24'd7781698, 24'd7662705, 24'd7687367, 24'd7850803, 24'd8120670, 24'd8443561, 24'd8755577, 24'd8994970, 24'd9114365, 24'd9090135, 24'd8927073, 24'd8657450, 24'd8334623, 24'd8022480, 24'd7782793, 24'd7662995, 24'd7686795, 24'd7849482, 24'd8118861, 24'd8441622, 24'd8753892, 24'd8993873, 24'd9114072, 24'd9090704, 24'd8928392, 24'd8659257, 24'd8336562, 24'd8024166, 24'd7783893, 
24'd7663291, 24'd7686228, 24'd7848165, 24'd8117055, 24'd8439684, 24'd8752205, 24'd8992771, 24'd9113774, 24'd9091268, 24'd8929707, 24'd8661063, 24'd8338501, 24'd8025854, 24'd7784996, 24'd7663592, 24'd7685666, 24'd7846852, 24'd8115250, 24'd8437745, 24'd8750515, 24'd8991665, 24'd9113471, 24'd9091828, 24'd8931018, 24'd8662867, 24'd8340440, 24'd8027545, 24'd7786104, 24'd7663897, 24'd7685109, 
24'd7845542, 24'd8113447, 24'd8435805, 24'd8748823, 24'd8990555, 24'd9113163, 24'd9092382, 24'd8932326, 24'd8664669, 24'd8342380, 24'd8029239, 24'd7787216, 24'd7664208, 24'd7684557, 24'd7844237, 24'd8111646, 24'd8433866, 24'd8747129, 24'd8989441, 24'd9112849, 24'd9092932, 24'd8933630, 24'd8666469, 24'd8344319, 24'd8030935, 24'd7788333, 24'd7664524, 24'd7684010, 24'd7842935, 24'd8109847, 
24'd8431926, 24'd8745431, 24'd8988322, 24'd9112531, 24'd9093476, 24'd8934930, 24'd8668267, 24'd8346260, 24'd8032633, 24'd7789453, 24'd7664845, 24'd7683468, 24'd7841637, 24'd8108050, 24'd8429985, 24'd8743732, 24'd8987200, 24'd9112207, 24'd9094016, 24'd8936226, 24'd8670063, 24'd8348200, 24'd8034334, 24'd7790578, 24'd7665171, 24'd7682931, 24'd7840343, 24'd8106255, 24'd8428045, 24'd8742029, 
24'd8986073, 24'd9111879, 24'd9094551, 24'd8937518, 24'd8671857, 24'd8350141, 24'd8036038, 24'd7791707, 24'd7665502, 24'd7682399, 24'd7839052, 24'd8104462, 24'd8426104, 24'd8740325, 24'd8984942, 24'd9111545, 24'd9095081, 24'd8938806, 24'd8673649, 24'd8352082, 24'd8037743, 24'd7792840, 24'd7665839, 24'd7681871, 24'd7837766, 24'd8102671, 24'd8424163, 24'd8738618, 24'd8983806, 24'd9111206, 
24'd9095605, 24'd8940091, 24'd8675439, 24'd8354023, 24'd8039452, 24'd7793978, 24'd7666180, 24'd7681349, 24'd7836483, 24'd8100882, 24'd8422221, 24'd8736908, 24'd8982667, 24'd9110863, 24'd9096125, 24'd8941371, 24'd8677227, 24'd8355965, 24'd8041163, 24'd7795119, 24'd7666526, 24'd7680832, 24'd7835205, 24'd8099095, 24'd8420279, 24'd8735196, 24'd8981523, 24'd9110514, 24'd9096640, 24'd8942648, 
24'd8679013, 24'd8357906, 24'd8042876, 24'd7796265, 24'd7666878, 24'd7680319, 24'd7833930, 24'd8097310, 24'd8418338, 24'd8733482, 24'd8980376, 24'd9110160, 24'd9097150, 24'd8943921, 24'd8680797, 24'd8359848, 24'd8044592, 24'd7797415, 24'd7667234, 24'd7679812, 24'd7832659, 24'd8095527, 24'd8416395, 24'd8731765, 24'd8979224, 24'd9109801, 24'd9097655, 24'd8945190, 24'd8682579, 24'd8361791, 
24'd8046310, 24'd7798569, 24'd7667596, 24'd7679309, 24'd7831392, 24'd8093746, 24'd8414453, 24'd8730045, 24'd8978068, 24'd9109437, 24'd9098155, 24'd8946455, 24'd8684358, 24'd8363733, 24'd8048030, 24'd7799727, 24'd7667962, 24'd7678812, 24'd7830129, 24'd8091967, 24'd8412511, 24'd8728324, 24'd8976907, 24'd9109068, 24'd9098650, 24'd8947716, 24'd8686136, 24'd8365676, 24'd8049753, 24'd7800889, 
24'd7668334, 24'd7678319, 24'd7828869, 24'd8090191, 24'd8410568, 24'd8726600, 24'd8975743, 24'd9108693, 24'd9099140, 24'd8948974, 24'd8687912, 24'd8367618, 24'd8051478, 24'd7802056, 24'd7668711, 24'd7677832, 24'd7827614, 24'd8088416, 24'd8408625, 24'd8724873, 24'd8974575, 24'd9108314, 24'd9099625, 24'd8950227, 24'd8689686, 24'd8369561, 24'd8053206, 24'd7803226, 24'd7669092, 24'd7677349, 
24'd7826363, 24'd8086643, 24'd8406682, 24'd8723144, 24'd8973402, 24'd9107930, 24'd9100105, 24'd8951477, 24'd8691457, 24'd8371504, 24'd8054936, 24'd7804401, 24'd7669479, 24'd7676872, 24'd7825115, 24'd8084873, 24'd8404739, 24'd8721413, 24'd8972225, 24'd9107541, 24'd9100580, 24'd8952722, 24'd8693226, 24'd8373447, 24'd8056668, 24'd7805579, 24'd7669871, 24'd7676399, 24'd7823872, 24'd8083105, 
24'd8402796, 24'd8719680, 24'd8971045, 24'd9107146, 24'd9101051, 24'd8953964, 24'd8694994, 24'd8375390, 24'd8058403, 24'd7806762, 24'd7670268, 24'd7675931, 24'd7822632, 24'd8081339, 24'd8400853, 24'd8717944, 24'd8969860, 24'd9106747, 24'd9101516, 24'd8955201, 24'd8696759, 24'd8377334, 24'd8060140, 24'd7807949, 24'd7670670, 24'd7675469, 24'd7821397, 24'd8079575, 24'd8398910, 24'd8716206, 
24'd8968671, 24'd9106343, 24'd9101976, 24'd8956435, 24'd8698522, 24'd8379277, 24'd8061879, 24'd7809140, 24'd7671077, 24'd7675011, 24'd7820165, 24'd8077813, 24'd8396966, 24'd8714465, 24'd8967478, 24'd9105933, 24'd9102431, 24'd8957664, 24'd8700282, 24'd8381221, 24'd8063621, 24'd7810335, 24'd7671488, 24'd7674558, 24'd7818937, 24'd8076053, 24'd8395023, 24'd8712723, 24'd8966281, 24'd9105519, 
24'd9102881, 24'd8958890, 24'd8702041, 24'd8383164, 24'd8065364, 24'd7811534, 24'd7671905, 24'd7674111, 24'd7817714, 24'd8074296, 24'd8393079, 24'd8710978, 24'd8965080, 24'd9105099, 24'd9103326, 24'd8960111, 24'd8703797, 24'd8385108, 24'd8067111, 24'd7812737, 24'd7672327, 24'd7673668, 24'd7816494, 24'd8072540, 24'd8391136, 24'd8709231, 24'd8963875, 24'd9104675, 24'd9103766, 24'd8961329, 
24'd8705551, 24'd8387051, 24'd8068859, 24'd7813944, 24'd7672755, 24'd7673231, 24'd7815279, 24'd8070787, 24'd8389192, 24'd8707481, 24'd8962666, 24'd9104245, 24'd9104201, 24'd8962543, 24'd8707303, 24'd8388995, 24'd8070610, 24'd7815155, 24'd7673187, 24'd7672798, 24'd7814067, 24'd8069037, 24'd8387248, 24'd8705729, 24'd8961452, 24'd9103811, 24'd9104631, 24'd8963752, 24'd8709053, 24'd8390938, 
24'd8072362, 24'd7816371, 24'd7673624, 24'd7672371, 24'd7812860, 24'd8067288, 24'd8385305, 24'd8703975, 24'd8960235, 24'd9103371, 24'd9105056, 24'd8964958, 24'd8710801, 24'd8392882, 24'd8074117, 24'd7817590, 24'd7674066, 24'd7671948, 24'd7811656, 24'd8065542, 24'd8383361, 24'd8702219, 24'd8959014, 24'd9102926, 24'd9105476, 24'd8966159, 24'd8712546, 24'd8394825, 24'd8075875, 24'd7818813, 
24'd7674513, 24'd7671531, 24'd7810457, 24'd8063798, 24'd8381418, 24'd8700461, 24'd8957789, 24'd9102477, 24'd9105891, 24'd8967357, 24'd8714289, 24'd8396769, 24'd8077634, 24'd7820040, 24'd7674965, 24'd7671118, 24'd7809261, 24'd8062056, 24'd8379474, 24'd8698700, 24'd8956560, 24'd9102022, 24'd9106301, 24'd8968550, 24'd8716029, 24'd8398712, 24'd8079396, 24'd7821271, 24'd7675422, 24'd7670711, 
24'd7808070, 24'd8060316, 24'd8377531, 24'd8696938, 24'd8955326, 24'd9101563, 24'd9106706, 24'd8969739, 24'd8717768, 24'd8400656, 24'd8081159, 24'd7822507, 24'd7675884, 24'd7670308, 24'd7806883, 24'd8058579, 24'd8375588, 24'd8695173, 24'd8954089, 24'd9101098, 24'd9107106, 24'd8970925, 24'd8719504, 24'd8402599, 24'd8082925, 24'd7823746, 24'd7676351, 24'd7669911, 24'd7805699, 24'd8056844, 
24'd8373644, 24'd8693406, 24'd8952848, 24'd9100628, 24'd9107501, 24'd8972106, 24'd8721237, 24'd8404542, 24'd8084693, 24'd7824989, 24'd7676823, 24'd7669519, 24'd7804520, 24'd8055112, 24'd8371701, 24'd8691637, 24'd8951603, 24'd9100154, 24'd9107891, 24'd8973283, 24'd8722969, 24'd8406485, 24'd8086464, 24'd7826236, 24'd7677300, 24'd7669131, 24'd7803345, 24'd8053381, 24'd8369758, 24'd8689865, 
24'd8950354, 24'd9099674, 24'd9108275, 24'd8974456, 24'd8724698, 24'd8408428, 24'd8088236, 24'd7827487, 24'd7677782, 24'd7668749, 24'd7802174, 24'd8051654, 24'd8367815, 24'd8688092, 24'd8949101, 24'd9099190, 24'd9108655, 24'd8975625, 24'd8726424, 24'd8410371, 24'd8090010, 24'd7828742, 24'd7678270, 24'd7668372, 24'd7801007, 24'd8049928, 24'd8365873, 24'd8686317, 24'd8947844, 24'd9098700, 
24'd9109030, 24'd8976789, 24'd8728149, 24'd8412314, 24'd8091787, 24'd7830001, 24'd7678762, 24'd7668000, 24'd7799845, 24'd8048205, 24'd8363930, 24'd8684539, 24'd8946583, 24'd9098206, 24'd9109399, 24'd8977950, 24'd8729871, 24'd8414256, 24'd8093566, 24'd7831263, 24'd7679259, 24'd7667633, 24'd7798686, 24'd8046484, 24'd8361988, 24'd8682759, 24'd8945319, 24'd9097706, 24'd9109764, 24'd8979106, 
24'd8731590, 24'd8416198, 24'd8095346, 24'd7832530, 24'd7679761, 24'd7667271, 24'd7797532, 24'd8044766, 24'd8360046, 24'd8680978, 24'd8944050, 24'd9097202, 24'd9110124, 24'd8980259, 24'd8733307, 24'd8418140, 24'd8097129, 24'd7833801, 24'd7680268, 24'd7666914, 24'd7796382, 24'd8043050, 24'd8358104, 24'd8679194, 24'd8942778, 24'd9096692, 24'd9110478, 24'd8981407, 24'd8735022, 24'd8420082, 
24'd8098914, 24'd7835075, 24'd7680779, 24'd7666562, 24'd7795235, 24'd8041336, 24'd8356162, 24'd8677408, 24'd8941501, 24'd9096178, 24'd9110827, 24'd8982551, 24'd8736734, 24'd8422024, 24'd8100701, 24'd7836353, 24'd7681296, 24'd7666215, 24'd7794093, 24'd8039625, 24'd8354220, 24'd8675620, 24'd8940221, 24'd9095658, 24'd9111172, 24'd8983691, 24'd8738444, 24'd8423965, 24'd8102489, 24'd7837636, 
24'd7681818, 24'd7665873, 24'd7792956, 24'd8037917, 24'd8352279, 24'd8673830, 24'd8938937, 24'd9095134, 24'd9111511, 24'd8984827, 24'd8740152, 24'd8425907, 24'd8104280, 24'd7838922, 24'd7682345, 24'd7665536, 24'd7791822, 24'd8036211, 24'd8350338, 24'd8672039, 24'd8937649, 24'd9094605, 24'd9111845, 24'd8985958, 24'd8741857, 24'd8427848, 24'd8106073, 24'd7840212, 24'd7682877, 24'd7665205, 
24'd7790693, 24'd8034507, 24'd8348397, 24'd8670245, 24'd8936357, 24'd9094071, 24'd9112174, 24'd8987085, 24'd8743559, 24'd8429788, 24'd8107868, 24'd7841505, 24'd7683413, 24'd7664878, 24'd7789567, 24'd8032806, 24'd8346457, 24'd8668449, 24'd8935061, 24'd9093531, 24'd9112498, 24'd8988209, 24'd8745259, 24'd8431729, 24'd8109665, 24'd7842803, 24'd7683955, 24'd7664557, 24'd7788446, 24'd8031107, 
24'd8344516, 24'd8666651, 24'd8933762, 24'd9092987, 24'd9112817, 24'd8989328, 24'd8746956, 24'd8433669, 24'd8111463, 24'd7844104, 24'd7684502, 24'd7664240, 24'd7787330, 24'd8029411, 24'd8342576, 24'd8664851, 24'd8932458, 24'd9092438, 24'd9113131, 24'd8990442, 24'd8748651, 24'd8435608, 24'd8113264, 24'd7845410, 24'd7685053, 24'd7663929, 24'd7786217, 24'd8027717, 24'd8340637, 24'd8663050, 
24'd8931151, 24'd9091884, 24'd9113440, 24'd8991553, 24'd8750344, 24'd8437548, 24'd8115067, 24'd7846719, 24'd7685610, 24'd7663622, 24'd7785109, 24'd8026026, 24'd8338698, 24'd8661246, 24'd8929840, 24'd9091325, 24'd9113744, 24'd8992659, 24'd8752034, 24'd8439487, 24'd8116871, 24'd7848032, 24'd7686171, 24'd7663321, 24'd7784004, 24'd8024337, 24'd8336759, 24'd8659441, 24'd8928526, 24'd9090761, 
24'd9114042, 24'd8993761, 24'd8753721, 24'd8441426, 24'd8118678, 24'd7849348, 24'd7686737, 24'd7663025, 24'd7782904, 24'd8022651, 24'd8334820, 24'd8657633, 24'd8927207, 24'd9090193, 24'd9114336, 24'd8994859, 24'd8755406, 24'd8443364, 24'd8120486, 24'd7850669, 24'd7687309, 24'd7662734, 24'd7781809, 24'd8020968, 24'd8332882, 24'd8655824, 24'd8925885, 24'd9089619, 24'd9114624, 24'd8995952, 
24'd8757088, 24'd8445302, 24'd8122296, 24'd7851993, 24'd7687885, 24'd7662448, 24'd7780717, 24'd8019287, 24'd8330944, 24'd8654013, 24'd8924559, 24'd9089040, 24'd9114908, 24'd8997042, 24'd8758768, 24'd8447240, 24'd8124108, 24'd7853321, 24'd7688466, 24'd7662167, 24'd7779630, 24'd8017609, 24'd8329007, 24'd8652200, 24'd8923229, 24'd9088457, 24'd9115186, 24'd8998127, 24'd8760445, 24'd8449177, 
24'd8125922, 24'd7854653, 24'd7689052, 24'd7661892, 24'd7778547, 24'd8015933, 24'd8327070, 24'd8650385, 24'd8921895, 24'd9087868, 24'd9115459, 24'd8999208, 24'd8762119, 24'd8451113, 24'd8127738, 24'd7855988, 24'd7689643, 24'd7661621, 24'd7777469, 24'd8014260, 24'd8325133, 24'd8648568, 24'd8920558, 24'd9087275, 24'd9115727, 24'd9000284, 24'd8763791, 24'd8453050, 24'd8129556, 24'd7857327, 
24'd7690238, 24'd7661355, 24'd7776394, 24'd8012589, 24'd8323197, 24'd8646750, 24'd8919217, 24'd9086677, 24'd9115990, 24'd9001356, 24'd8765460, 24'd8454986, 24'd8131375, 24'd7858670, 24'd7690839, 24'd7661095, 24'd7775324, 24'd8010921, 24'd8321262, 24'd8644930, 24'd8917872, 24'd9086074, 24'd9116248, 24'd9002424, 24'd8767127, 24'd8456921, 24'd8133196, 24'd7860017, 24'd7691445, 24'd7660840, 
24'd7774259, 24'd8009256, 24'd8319327, 24'd8643108, 24'd8916523, 24'd9085466, 24'd9116501, 24'd9003488, 24'd8768791, 24'd8458856, 24'd8135019, 24'd7861367, 24'd7692055, 24'd7660589, 24'd7773197, 24'd8007594, 24'd8317392, 24'd8641284, 24'd8915171, 24'd9084853, 24'd9116749, 24'd9004547, 24'd8770452, 24'd8460790, 24'd8136844, 24'd7862721, 24'd7692670, 24'd7660344, 24'd7772140, 24'd8005934, 
24'd8315458, 24'd8639458, 24'd8913815, 24'd9084235, 24'd9116991, 24'd9005602, 24'd8772110, 24'd8462724, 24'd8138671, 24'd7864079, 24'd7693291, 24'd7660104, 24'd7771087, 24'd8004276, 24'd8313524, 24'd8637631, 24'd8912456, 24'd9083612, 24'd9117229, 24'd9006652, 24'd8773766, 24'd8464658, 24'd8140499, 24'd7865440, 24'd7693916, 24'd7659869, 24'd7770039, 24'd8002622, 24'd8311591, 24'd8635801, 
24'd8911093, 24'd9082985, 24'd9117461, 24'd9007699, 24'd8775419, 24'd8466590, 24'd8142329, 24'd7866805, 24'd7694546, 24'd7659640, 24'd7768995, 24'd8000970, 24'd8309658, 24'd8633970, 24'd8909726, 24'd9082352, 24'd9117688, 24'd9008741, 24'd8777070, 24'd8468523, 24'd8144161, 24'd7868174, 24'd7695181, 24'd7659415, 24'd7767955, 24'd7999321, 24'd8307726, 24'd8632138, 24'd8908355, 24'd9081715, 
24'd9117911, 24'd9009778, 24'd8778717, 24'd8470454, 24'd8145994, 24'd7869547, 24'd7695820, 24'd7659195, 24'd7766920, 24'd7997675, 24'd8305795, 24'd8630303, 24'd8906981, 24'd9081073, 24'd9118128, 24'd9010812, 24'd8780362, 24'd8472386, 24'd8147829, 24'd7870923, 24'd7696465, 24'd7658981, 24'd7765888, 24'd7996031, 24'd8303864, 24'd8628467, 24'd8905603, 24'd9080426, 24'd9118340, 24'd9011840, 
24'd8782005, 24'd8474316, 24'd8149666, 24'd7872302, 24'd7697114, 24'd7658771, 24'd7764862, 24'd7994390, 24'd8301934, 24'd8626630, 24'd8904222, 24'd9079774, 24'd9118546, 24'd9012865, 24'd8783644, 24'd8476246, 24'd8151505, 24'd7873686, 24'd7697768, 24'd7658567, 24'd7763839, 24'd7992752, 24'd8300004, 24'd8624790, 24'd8902836, 24'd9079118, 24'd9118748, 24'd9013885, 24'd8785281, 24'd8478176, 
24'd8153345, 24'd7875072, 24'd7698428, 24'd7658368, 24'd7762821, 24'd7991117, 24'd8298075, 24'd8622949, 24'd8901448, 24'd9078456, 24'd9118945, 24'd9014901, 24'd8786915, 24'd8480104, 24'd8155187, 24'd7876463, 24'd7699091, 24'd7658174, 24'd7761808, 24'd7989484, 24'd8296147, 24'd8621107, 24'd8900056, 24'd9077790, 24'd9119136, 24'd9015912, 24'd8788546, 24'd8482032, 24'd8157030, 24'd7877857, 
24'd7699760, 24'd7657985, 24'd7760799, 24'd7987855, 24'd8294219, 24'd8619262, 24'd8898660, 24'd9077119, 24'd9119322, 24'd9016919, 24'd8790174, 24'd8483960, 24'd8158875, 24'd7879255, 24'd7700434, 24'd7657801, 24'd7759794, 24'd7986228, 24'd8292292, 24'd8617416, 24'd8897260, 24'd9076443, 24'd9119504, 24'd9017922, 24'd8791800, 24'd8485887, 24'd8160722, 24'd7880656, 24'd7701112, 24'd7657623, 
24'd7758794, 24'd7984604, 24'd8290365, 24'd8615569, 24'd8895857, 24'd9075762, 24'd9119680, 24'd9018920, 24'd8793422, 24'd8487813, 24'd8162571, 24'd7882061, 24'd7701795, 24'd7657449, 24'd7757798, 24'd7982982, 24'd8288440, 24'd8613720, 24'd8894451, 24'd9075076, 24'd9119851, 24'd9019914, 24'd8795042, 24'd8489738, 24'd8164420, 24'd7883469, 24'd7702484, 24'd7657281, 24'd7756806, 24'd7981364, 
24'd8286515, 24'd8611869, 24'd8893041, 24'd9074386, 24'd9120017, 24'd9020903, 24'd8796659, 24'd8491663, 24'd8166272, 24'd7884881, 24'd7703176, 24'd7657118, 24'd7755819, 24'd7979748, 24'd8284590, 24'd8610017, 24'd8891627, 24'd9073690, 24'd9120177, 24'd9021888, 24'd8798273, 24'd8493587, 24'd8168125, 24'd7886296, 24'd7703874, 24'd7656959, 24'd7754836, 24'd7978136, 24'd8282667, 24'd8608163, 
24'd8890210, 24'd9072990, 24'd9120333, 24'd9022868, 24'd8799885, 24'd8495510, 24'd8169980, 24'd7887715, 24'd7704577, 24'd7656806, 24'd7753858, 24'd7976526, 24'd8280744, 24'd8606308, 24'd8888789, 24'd9072285, 24'd9120483, 24'd9023844, 24'd8801493, 24'd8497432, 24'd8171836, 24'd7889138, 24'd7705284, 24'd7656658, 24'd7752885, 24'd7974919, 24'd8278822, 24'd8604451, 24'd8887365, 24'd9071576, 
24'd9120629, 24'd9024816, 24'd8803098, 24'd8499354, 24'd8173693, 24'd7890564, 24'd7705996, 24'd7656516, 24'd7751915, 24'd7973315, 24'd8276900, 24'd8602592, 24'd8885937, 24'd9070861, 24'd9120769, 24'd9025783, 24'd8804701, 24'd8501275, 24'd8175552, 24'd7891993, 24'd7706713, 24'd7656378, 24'd7750950, 24'd7971714, 24'd8274980, 24'd8600732, 24'd8884506, 24'd9070142, 24'd9120904, 24'd9026745, 
24'd8806301, 24'd8503195, 24'd8177413, 24'd7893426, 24'd7707434, 24'd7656246, 24'd7749990, 24'd7970116, 24'd8273060, 24'd8598871, 24'd8883071, 24'd9069418, 24'd9121034, 24'd9027703, 24'd8807897, 24'd8505115, 24'd8179275, 24'd7894862, 24'd7708161, 24'd7656118, 24'd7749034, 24'd7968520, 24'd8271141, 24'd8597008, 24'd8881633, 24'd9068689, 24'd9121158, 24'd9028657, 24'd8809491, 24'd8507033, 
24'd8181139, 24'd7896302, 24'd7708892, 24'd7655996, 24'd7748083, 24'd7966928, 24'd8269223, 24'd8595144, 24'd8880192, 24'd9067956, 24'd9121278, 24'd9029606, 24'd8811082, 24'd8508951, 24'd8183004, 24'd7897746, 24'd7709628, 24'd7655879, 24'd7747136, 24'd7965339, 24'd8267306, 24'd8593278, 24'd8878747, 24'd9067217, 24'd9121393, 24'd9030551, 24'd8812670, 24'd8510868, 24'd8184870, 24'd7899192, 
24'd7710369, 24'd7655767, 24'd7746193, 24'd7963752, 24'd8265389, 24'd8591411, 24'd8877298, 24'd9066474, 24'd9121502, 24'd9031491, 24'd8814255, 24'd8512784, 24'd8186738, 24'd7900642, 24'd7711114, 24'd7655660, 24'd7745256, 24'd7962169, 24'd8263474, 24'd8589542, 24'd8875846, 24'd9065726, 24'd9121606, 24'd9032427, 24'd8815837, 24'd8514699, 24'd8188608, 24'd7902096, 24'd7711864, 24'd7655559, 
24'd7744322, 24'd7960588, 24'd8261559, 24'd8587672, 24'd8874391, 24'd9064974, 24'd9121705, 24'd9033358, 24'd8817416, 24'd8516613, 24'd8190478, 24'd7903553, 24'd7712619, 24'd7655462, 24'd7743393, 24'd7959011, 24'd8259645, 24'd8585801, 24'd8872932, 24'd9064217, 24'd9121799, 24'd9034284, 24'd8818992, 24'd8518526, 24'd8192350, 24'd7905014, 24'd7713379, 24'd7655371, 24'd7742469, 24'd7957437, 
24'd8257732, 24'd8583928, 24'd8871470, 24'd9063454, 24'd9121888, 24'd9035207, 24'd8820564, 24'd8520439, 24'd8194224, 24'd7906477, 24'd7714143, 24'd7655285, 24'd7741549, 24'd7955865, 24'd8255820, 24'd8582054, 24'd8870005, 24'd9062688, 24'd9121972, 24'd9036124, 24'd8822134, 24'd8522350, 24'd8196099, 24'd7907945, 24'd7714912, 24'd7655203, 24'd7740634, 24'd7954297, 24'd8253909, 24'd8580178, 
24'd8868536, 24'd9061916, 24'd9122050, 24'd9037037, 24'd8823701, 24'd8524261, 24'd8197975, 24'd7909415, 24'd7715686, 24'd7655128, 24'd7739723, 24'd7952732, 24'd8251999, 24'd8578301, 24'd8867063, 24'd9061140, 24'd9122123, 24'd9037946, 24'd8825265, 24'd8526170, 24'd8199853, 24'd7910889, 24'd7716465, 24'd7655057, 24'd7738817, 24'd7951169, 24'd8250090, 24'd8576423, 24'd8865588, 24'd9060359, 
24'd9122192, 24'd9038850, 24'd8826826, 24'd8528079, 24'd8201731, 24'd7912366, 24'd7717248, 24'd7654991, 24'd7737915, 24'd7949610, 24'd8248182, 24'd8574544, 24'd8864109, 24'd9059573, 24'd9122255, 24'd9039749, 24'd8828383, 24'd8529987, 24'd8203612, 24'd7913847, 24'd7718036, 24'd7654931, 24'd7737018, 24'd7948054, 24'd8246275, 24'd8572663, 24'd8862627, 24'd9058783, 24'd9122313, 24'd9040644, 
24'd8829938, 24'd8531893, 24'd8205493, 24'd7915331, 24'd7718829, 24'd7654875, 24'd7736126, 24'd7946501, 24'd8244369, 24'd8570781, 24'd8861141, 24'd9057988, 24'd9122366, 24'd9041534, 24'd8831489, 24'd8533799, 24'd8207376, 24'd7916818, 24'd7719626, 24'd7654825, 24'd7735238, 24'd7944951, 24'd8242463, 24'd8568897, 24'd8859652, 24'd9057188, 24'd9122413, 24'd9042420, 24'd8833038, 24'd8535704, 
24'd8209260, 24'd7918309, 24'd7720429, 24'd7654780, 24'd7734354, 24'd7943404, 24'd8240559, 24'd8567013, 24'd8858160, 24'd9056384, 24'd9122456, 24'd9043301, 24'd8834583, 24'd8537607, 24'd8211145, 24'd7919802, 24'd7721235, 24'd7654740, 24'd7733476, 24'd7941861, 24'd8238656, 24'd8565127, 24'd8856664, 24'd9055575, 24'd9122493, 24'd9044177, 24'd8836125, 24'd8539510, 24'd8213032, 24'd7921300, 
24'd7722047, 24'd7654705, 24'd7732601, 24'd7940320, 24'd8236754, 24'd8563240, 24'd8855166, 24'd9054761, 24'd9122525, 24'd9045049, 24'd8837664, 24'd8541412, 24'd8214920, 24'd7922800, 24'd7722863, 24'd7654676, 24'd7731732, 24'd7938783, 24'd8234853, 24'd8561351, 24'd8853664, 24'd9053942, 24'd9122552, 24'd9045916, 24'd8839200, 24'd8543312, 24'd8216809, 24'd7924304, 24'd7723684, 24'd7654651, 
24'd7730867, 24'd7937248, 24'd8232953, 24'd8559462, 24'd8852158, 24'd9053119, 24'd9122574, 24'd9046779, 24'd8840732, 24'd8545211, 24'd8218699, 24'd7925811, 24'd7724509, 24'd7654632, 24'd7730007, 24'd7935717, 24'd8231054, 24'd8557571, 24'd8850650, 24'd9052291, 24'd9122591, 24'd9047637, 24'd8842262, 24'd8547110, 24'd8220590, 24'd7927321, 24'd7725339, 24'd7654617, 24'd7729151, 24'd7934189, 
24'd8229157, 24'd8555679, 24'd8849138, 24'd9051459, 24'd9122603, 24'd9048490, 24'd8843788, 24'd8549007, 24'd8222483, 24'd7928834, 24'd7726174, 24'd7654608, 24'd7728300, 24'd7932665, 24'd8227260, 24'd8553786, 24'd8847623, 24'd9050622, 24'd9122609, 24'd9049339, 24'd8845311, 24'd8550903, 24'd8224376, 24'd7930351, 24'd7727014, 24'd7654604, 24'd7727453, 24'd7931143, 24'd8225365, 24'd8551891, 
24'd8846105, 24'd9049780, 24'd9122611, 24'd9050183, 24'd8846831, 24'd8552798, 24'd8226271, 24'd7931871, 24'd7727858, 24'd7654606, 24'd7726611, 24'd7929625, 24'd8223470, 24'd8549996, 24'd8844583, 24'd9048934, 24'd9122607, 24'd9051023, 24'd8848348, 24'd8554692, 24'd8228167, 24'd7933394, 24'd7728706, 24'd7654612, 24'd7725774, 24'd7928110, 24'd8221577, 24'd8548099, 24'd8843058, 24'd9048083, 
24'd9122598, 24'd9051858, 24'd8849862, 24'd8556584, 24'd8230064, 24'd7934920, 24'd7729560, 24'd7654624, 24'd7724942, 24'd7926598, 24'd8219685, 24'd8546202, 24'd8841531, 24'd9047227, 24'd9122584, 24'd9052688, 24'd8851372, 24'd8558476, 24'd8231963, 24'd7936450, 24'd7730418, 24'd7654640, 24'd7724114, 24'd7925089, 24'd8217794, 24'd8544303, 24'd8840000, 24'd9046367, 24'd9122564, 24'd9053513, 
24'd8852879, 24'd8560366, 24'd8233862, 24'd7937982, 24'd7731280, 24'd7654662, 24'd7723290, 24'd7923584, 24'd8215905, 24'd8542403, 24'd8838465, 24'd9045502, 24'd9122540, 24'd9054334, 24'd8854383, 24'd8562255, 24'd8235762, 24'd7939518, 24'd7732147, 24'd7654689, 24'd7722472, 24'd7922082, 24'd8214016, 24'd8540502, 24'd8836928, 24'd9044632, 24'd9122511, 24'd9055151, 24'd8855883, 24'd8564143, 
24'd8237664, 24'd7941057, 24'd7733019, 24'd7654721, 24'd7721658, 24'd7920583, 24'd8212129, 24'd8538600, 24'd8835388, 24'd9043758, 24'd9122476, 24'd9055962, 24'd8857380, 24'd8566029, 24'd8239567, 24'd7942599, 24'd7733895, 24'd7654758, 24'd7720849, 24'd7919087, 24'd8210243, 24'd8536697, 24'd8833844, 24'd9042880, 24'd9122436, 24'd9056769, 24'd8858874, 24'd8567914, 24'd8241470, 24'd7944144, 
24'd7734776, 24'd7654801, 24'd7720044, 24'd7917595, 24'd8208358, 24'd8534793, 24'd8832297, 24'd9041996, 24'd9122391, 24'd9057571, 24'd8860365, 24'd8569798, 24'd8243375, 24'd7945692, 24'd7735662, 24'd7654848, 24'd7719244, 24'd7916106, 24'd8206475, 24'd8532888, 24'd8830747, 24'd9041109, 24'd9122341, 24'd9058369, 24'd8861852, 24'd8571681, 24'd8245280, 24'd7947244, 24'd7736552, 24'd7654901, 
24'd7718449, 24'd7914620, 24'd8204593, 24'd8530981, 24'd8829194, 24'd9040216, 24'd9122286, 24'd9059162, 24'd8863336, 24'd8573563, 24'd8247187, 24'd7948798, 24'd7737447, 24'd7654959, 24'd7717659, 24'd7913138, 24'd8202712, 24'd8529074, 24'd8827638, 24'd9039319, 24'd9122225, 24'd9059950, 24'd8864817, 24'd8575443, 24'd8249095, 24'd7950356, 24'd7738346, 24'd7655022, 24'd7716873, 24'd7911659, 
24'd8200832, 24'd8527166, 24'd8826079, 24'd9038418, 24'd9122160, 24'd9060733, 24'd8866294, 24'd8577322, 24'd8251003, 24'd7951916, 24'd7739250, 24'd7655090, 24'd7716092, 24'd7910183, 24'd8198954, 24'd8525257, 24'd8824517, 24'd9037512, 24'd9122089, 24'd9061512, 24'd8867768, 24'd8579199, 24'd8252913, 24'd7953480, 24'd7740158, 24'd7655163, 24'd7715316, 24'd7908711, 24'd8197077, 24'd8523347, 
24'd8822952, 24'd9036601, 24'd9122013, 24'd9062286, 24'd8869239, 24'd8581076, 24'd8254824, 24'd7955047, 24'd7741071, 24'd7655242, 24'd7714544, 24'd7907242, 24'd8195202, 24'd8521436, 24'd8821384, 24'd9035686, 24'd9121932, 24'd9063055, 24'd8870706, 24'd8582951, 24'd8256735, 24'd7956617, 24'd7741989, 24'd7655325, 24'd7713777, 24'd7905777, 24'd8193327, 24'd8519524, 24'd8819812, 24'd9034766, 
24'd9121846, 24'd9063820, 24'd8872170, 24'd8584824, 24'd8258647, 24'd7958190, 24'd7742911, 24'd7655414, 24'd7713015, 24'd7904314, 24'd8191455, 24'd8517611, 24'd8818238, 24'd9033842, 24'd9121755, 24'd9064579, 24'd8873630, 24'd8586696, 24'd8260561, 24'd7959765, 24'd7743837, 24'd7655508, 24'd7712257, 24'd7902856, 24'd8189583, 24'd8515697, 24'd8816661, 24'd9032913, 24'd9121658, 24'd9065335, 
24'd8875088, 24'd8588567, 24'd8262475, 24'd7961344, 24'd7744768, 24'd7655607, 24'd7711505, 24'd7901400, 24'd8187713, 24'd8513783, 24'd8815080, 24'd9031980, 24'd9121557, 24'd9066085, 24'd8876541, 24'd8590436, 24'd8264390, 24'd7962926, 24'd7745704, 24'd7655711, 24'd7710757, 24'd7899948, 24'd8185844, 24'd8511867, 24'd8813497, 24'd9031042, 24'd9121450, 24'd9066830, 24'd8877991, 24'd8592304, 
24'd8266306, 24'd7964511, 24'd7746644, 24'd7655820, 24'd7710014, 24'd7898500, 24'd8183977, 24'd8509951, 24'd8811911, 24'd9030100, 24'd9121338, 24'd9067571, 24'd8879438, 24'd8594171, 24'd8268223, 24'd7966099, 24'd7747588, 24'd7655934, 24'd7709275, 24'd7897055, 24'd8182111, 24'd8508033, 24'd8810321, 24'd9029153, 24'd9121221, 24'd9068307, 24'd8880882, 24'd8596036, 24'd8270141, 24'd7967690, 
24'd7748537, 24'd7656054, 24'd7708542, 24'd7895613, 24'd8180247, 24'd8506115, 24'd8808729, 24'd9028201, 24'd9121099, 24'd9069039, 24'd8882322, 24'd8597900, 24'd8272059, 24'd7969283, 24'd7749491, 24'd7656179, 24'd7707813, 24'd7894175, 24'd8178384, 24'd8504196, 24'd8807134, 24'd9027246, 24'd9120972, 24'd9069765, 24'd8883758, 24'd8599762, 24'd8273978, 24'd7970880, 24'd7750449, 24'd7656308, 
24'd7707089, 24'd7892740, 24'd8176523, 24'd8502277, 24'd8805536, 24'd9026285, 24'd9120840, 24'd9070487, 24'd8885191, 24'd8601622, 24'd8275899, 24'd7972480, 24'd7751411, 24'd7656443, 24'd7706369, 24'd7891309, 24'd8174663, 24'd8500356, 24'd8803935, 24'd9025321, 24'd9120702, 24'd9071204, 24'd8886621, 24'd8603482, 24'd8277819, 24'd7974082, 24'd7752378, 24'd7656583, 24'd7705655, 24'd7889881, 
24'd8172804, 24'd8498435, 24'd8802331, 24'd9024351, 24'd9120560, 24'd9071916, 24'd8888047, 24'd8605339, 24'd8279741, 24'd7975687, 24'd7753350, 24'd7656729, 24'd7704945, 24'd7888457, 24'd8170947, 24'd8496513, 24'd8800724, 24'd9023378, 24'd9120412, 24'd9072623, 24'd8889469, 24'd8607195, 24'd8281664, 24'd7977296, 24'd7754326, 24'd7656879, 24'd7704240, 24'd7887036, 24'd8169092, 24'd8494590, 
24'd8799114, 24'd9022400, 24'd9120259, 24'd9073326, 24'd8890888, 24'd8609050, 24'd8283587, 24'd7978907, 24'd7755306, 24'd7657034, 24'd7703540, 24'd7885619, 24'd8167238, 24'd8492666, 24'd8797501, 24'd9021417, 24'd9120101, 24'd9074024, 24'd8892304, 24'd8610903, 24'd8285511, 24'd7980521, 24'd7756291, 24'd7657195, 24'd7702844, 24'd7884205, 24'd8165386, 24'd8490742, 24'd8795886, 24'd9020430, 
24'd9119938, 24'd9074717, 24'd8893716, 24'd8612755, 24'd8287435, 24'd7982138, 24'd7757280, 24'd7657361, 24'd7702154, 24'd7882795, 24'd8163535, 24'd8488817, 24'd8794268, 24'd9019439, 24'd9119770, 24'd9075405, 24'd8895124, 24'd8614605, 24'd8289361, 24'd7983758, 24'd7758274, 24'd7657532, 24'd7701468, 24'd7881388, 24'd8161686, 24'd8486891, 24'd8792646, 24'd9018443, 24'd9119596, 24'd9076088, 
24'd8896529, 24'd8616453, 24'd8291287, 24'd7985380, 24'd7759272, 24'd7657708, 24'd7700787, 24'd7879985, 24'd8159838, 24'd8484965, 24'd8791022, 24'd9017443, 24'd9119418, 24'd9076767, 24'd8897930, 24'd8618300, 24'd8293214, 24'd7987006, 24'd7760274, 24'd7657889, 24'd7700111, 24'd7878585, 24'd8157992, 24'd8483038, 24'd8789395, 24'd9016438, 24'd9119234, 24'd9077440, 24'd8899328, 24'd8620145, 
24'd8295141, 24'd7988634, 24'd7761281, 24'd7658075, 24'd7699440, 24'd7877190, 24'd8156148, 24'd8481110, 24'd8787766, 24'd9015429, 24'd9119045, 24'd9078109, 24'd8900722, 24'd8621988, 24'd8297069, 24'd7990265, 24'd7762292, 24'd7658266, 24'd7698773, 24'd7875797, 24'd8154305, 24'd8479182, 24'd8786133, 24'd9014415, 24'd9118851, 24'd9078773, 24'd8902113, 24'd8623830, 24'd8298998, 24'd7991899, 
24'd7763308, 24'd7658463, 24'd7698112, 24'd7874408, 24'd8152464, 24'd8477253, 24'd8784498, 24'd9013398, 24'd9118652, 24'd9079432, 24'd8903500, 24'd8625671, 24'd8300927, 24'd7993536, 24'd7764328, 24'd7658664, 24'd7697455, 24'd7873023, 24'd8150625, 24'd8475323, 24'd8782860, 24'd9012375, 24'd9118448, 24'd9080087, 24'd8904883, 24'd8627509, 24'd8302857, 24'd7995175, 24'd7765352, 24'd7658871, 
24'd7696803, 24'd7871642, 24'd8148787, 24'd8473393, 24'd8781219, 24'd9011349, 24'd9118239, 24'd9080736, 24'd8906263, 24'd8629346, 24'd8304788, 24'd7996817, 24'd7766381, 24'd7659083, 24'd7696156, 24'd7870264, 24'd8146951, 24'd8471462, 24'd8779576, 24'd9010318, 24'd9118024, 24'd9081381, 24'd8907639, 24'd8631181, 24'd8306719, 24'd7998462, 24'd7767414, 24'd7659300, 24'd7695514, 24'd7868890, 
24'd8145117, 24'd8469530, 24'd8777929, 24'd9009282, 24'd9117805, 24'd9082021, 24'd8909011, 24'd8633015, 24'd8308651, 24'd8000110, 24'd7768452, 24'd7659522, 24'd7694876, 24'd7867519, 24'd8143284, 24'd8467598, 24'd8776280, 24'd9008243, 24'd9117580, 24'd9082656, 24'd8910380, 24'd8634847, 24'd8310583, 24'd8001760, 24'd7769494, 24'd7659749, 24'd7694244, 24'd7866152, 24'd8141453, 24'd8465666, 
24'd8774629, 24'd9007199, 24'd9117351, 24'd9083286, 24'd8911745, 24'd8636677, 24'd8312516, 24'd8003413, 24'd7770540, 24'd7659981, 24'd7693616, 24'd7864789, 24'd8139624, 24'd8463733, 24'd8772974, 24'd9006150, 24'd9117116, 24'd9083911, 24'd8913107, 24'd8638505, 24'd8314449, 24'd8005069, 24'd7771590, 24'd7660218, 24'd7692993, 24'd7863429, 24'd8137796, 24'd8461799, 24'd8771317, 24'd9005098, 
24'd9116876, 24'd9084531, 24'd8914465, 24'd8640332, 24'd8316383, 24'd8006728, 24'd7772645, 24'd7660461, 24'd7692375, 24'd7862073, 24'd8135971, 24'd8459865, 24'd8769657, 24'd9004041, 24'd9116631, 24'd9085147, 24'd8915819, 24'd8642156, 24'd8318317, 24'd8008389, 24'd7773705, 24'd7660709, 24'd7691762, 24'd7860721, 24'd8134147, 24'd8457930, 24'd8767995, 24'd9002979, 24'd9116381, 24'd9085757, 
24'd8917169, 24'd8643980, 24'd8320252, 24'd8010052, 24'd7774768, 24'd7660961, 24'd7691154, 24'd7859372, 24'd8132325, 24'd8455995, 24'd8766330, 24'd9001914, 24'd9116126, 24'd9086363, 24'd8918516, 24'd8645801, 24'd8322188, 24'd8011719, 24'd7775836, 24'd7661219, 24'd7690551, 24'd7858027, 24'd8130504, 24'd8454059, 24'd8764662, 24'd9000844, 24'd9115865, 24'd9086964, 24'd8919859, 24'd8647620, 
24'd8324124, 24'd8013388, 24'd7776908, 24'd7661482, 24'd7689953, 24'd7856686, 24'd8128686, 24'd8452123, 24'd8762991, 24'd8999769, 24'd9115600, 24'd9087560, 24'd8921198, 24'd8649438, 24'd8326060, 24'd8015060, 24'd7777984, 24'd7661750, 24'd7689359, 24'd7855349, 24'd8126869, 24'd8450187, 24'd8761318, 24'd8998691, 24'd9115329, 24'd9088151, 24'd8922534, 24'd8651254, 24'd8327997, 24'd8016734, 
24'd7779065, 24'd7662023, 24'd7688771, 24'd7854015, 24'd8125054, 24'd8448250, 24'd8759643, 24'd8997608, 24'd9115054, 24'd9088737, 24'd8923865, 24'd8653068, 24'd8329934, 24'd8018411, 24'd7780150, 24'd7662301, 24'd7688187, 24'd7852685, 24'd8123241, 24'd8446313, 24'd8757964, 24'd8996521, 24'd9114773, 24'd9089318, 24'd8925193, 24'd8654880, 24'd8331871, 24'd8020091, 24'd7781239, 24'd7662584, 
24'd7687608, 24'd7851359, 24'd8121430, 24'd8444375, 24'd8756284, 24'd8995430, 24'd9114487, 24'd9089894, 24'd8926518, 24'd8656690, 24'd8333809, 24'd8021773, 24'd7782332, 24'd7662873, 24'd7687035, 24'd7850037, 24'd8119621, 24'd8442437, 24'd8754600, 24'd8994334, 24'd9114196, 24'd9090465, 24'd8927838, 24'd8658498, 24'd8335748, 24'd8023458, 24'd7783430, 24'd7663166, 24'd7686466, 24'd7848718, 
24'd8117813, 24'd8440498, 24'd8752914, 24'd8993234, 24'd9113900, 24'd9091032, 24'd8929155, 24'd8660305, 24'd8337686, 24'd8025145, 24'd7784532, 24'd7663465, 24'd7685902, 24'd7847403, 24'd8116008, 24'd8438559, 24'd8751225, 24'd8992130, 24'd9113599, 24'd9091593, 24'd8930468, 24'd8662109, 24'd8339625, 24'd8026835, 24'd7785638, 24'd7663768, 24'd7685343, 24'd7846092, 24'd8114204, 24'd8436620, 
24'd8749534, 24'd8991022, 24'd9113293, 24'd9092150, 24'd8931777, 24'd8663912, 24'd8341565, 24'd8028527, 24'd7786749, 24'd7664077, 24'd7684789, 24'd7844785, 24'd8112402, 24'd8434680, 24'd8747841, 24'd8989909, 24'd9112982, 24'd9092702, 24'd8933082, 24'd8665713, 24'd8343504, 24'd8030222, 24'd7787863, 24'd7664391, 24'd7684240, 24'd7843481, 24'd8110603, 24'd8432741, 24'd8746145, 24'd8988793, 
24'd9112665, 24'd9093248, 24'd8934384, 24'd8667512, 24'd8345445, 24'd8031919, 24'd7788982, 24'd7664710, 24'd7683695, 24'd7842182, 24'd8108805, 24'd8430800, 24'd8744446, 24'd8987672, 24'd9112344, 24'd9093790, 24'd8935682, 24'd8669308, 24'd8347385, 24'd8033619, 24'd7790105, 24'd7665034, 24'd7683156, 24'd7840886, 24'd8107009, 24'd8428860, 24'd8742745, 24'd8986547, 24'd9112017, 24'd9094327, 
24'd8936976, 24'd8671103, 24'd8349326, 24'd8035322, 24'd7791232, 24'd7665363, 24'd7682622, 24'd7839594, 24'd8105215, 24'd8426919, 24'd8741041, 24'd8985417, 24'd9111686, 24'd9094859, 24'd8938266, 24'd8672896, 24'd8351267, 24'd8037027, 24'd7792364, 24'd7665697, 24'd7682092, 24'd7838306, 24'd8103423, 24'd8424978, 24'd8739335, 24'd8984284, 24'd9111349, 24'd9095386, 24'd8939552, 24'd8674687, 
24'd8353208, 24'd8038734, 24'd7793500, 24'd7666036, 24'd7681568, 24'd7837022, 24'd8101633, 24'd8423037, 24'd8737626, 24'd8983146, 24'd9111008, 24'd9095907, 24'd8940834, 24'd8676476, 24'd8355149, 24'd8040444, 24'd7794639, 24'd7666380, 24'd7681048, 24'd7835741, 24'd8099845, 24'd8421095, 24'd8735915, 24'd8982004, 24'd9110661, 24'd9096424, 24'd8942112, 24'd8678263, 24'd8357091, 24'd8042156, 
24'd7795783, 24'd7666729, 24'd7680534, 24'd7834465, 24'd8098060, 24'd8419153, 24'd8734202, 24'd8980858, 24'd9110309, 24'd9096937, 24'd8943387, 24'd8680048, 24'd8359033, 24'd8043871, 24'd7796931, 24'd7667084, 24'd7680024, 24'd7833192, 24'd8096276, 24'd8417211, 24'd8732486, 24'd8979708, 24'd9109952, 24'd9097444, 24'd8944658, 24'd8681830, 24'd8360975, 24'd8045588, 24'd7798084, 24'd7667443, 
24'd7679520, 24'd7831924, 24'd8094494, 24'd8415269, 24'd8730768, 24'd8978554, 24'd9109590, 24'd9097946, 24'd8945924, 24'd8683611, 24'd8362917, 24'd8047307, 24'd7799240, 24'd7667808, 24'd7679020, 24'd7830659, 24'd8092714, 24'd8413327, 24'd8729047, 24'd8977395, 24'd9109223, 24'd9098443, 24'd8947187, 24'd8685390, 24'd8364860, 24'd8049029, 24'd7800401, 24'd7668177, 24'd7678526, 24'd7829398, 
24'd8090937, 24'd8411384, 24'd8727324, 24'd8976233, 24'd9108851, 24'd9098935, 24'd8948446, 24'd8687166, 24'd8366802, 24'd8050753, 24'd7801565, 24'd7668552, 24'd7678036, 24'd7828141, 24'd8089161, 24'd8409441, 24'd8725599, 24'd8975066, 24'd9108474, 24'd9099422, 24'd8949701, 24'd8688941, 24'd8368745, 24'd8052480, 24'd7802734, 24'd7668931, 24'd7677551, 24'd7826888, 24'd8087388, 24'd8407499, 
24'd8723871, 24'd8973895, 24'd9108092, 24'd9099904, 24'd8950952, 24'd8690713, 24'd8370688, 24'd8054209, 24'd7803907, 24'd7669316, 24'd7677072, 24'd7825639, 24'd8085616, 24'd8405556, 24'd8722141, 24'd8972720, 24'd9107705, 24'd9100381, 24'd8952199, 24'd8692483, 24'd8372631, 24'd8055940, 24'd7805084, 24'd7669706, 24'd7676597, 24'd7824394, 24'd8083847, 24'd8403612, 24'd8720408, 24'd8971541, 
24'd9107313, 24'd9100854, 24'd8953443, 24'd8694252, 24'd8374574, 24'd8057674, 24'd7806265, 24'd7670100, 24'd7676127, 24'd7823152, 24'd8082080, 24'd8401669, 24'd8718673, 24'd8970358, 24'd9106915, 24'd9101321, 24'd8954682, 24'd8696018, 24'd8376517, 24'd8059410, 24'd7807450, 24'd7670500, 24'd7675662, 24'd7821915, 24'd8080315, 24'd8399726, 24'd8716936, 24'd8969171, 24'd9106513, 24'd9101783, 
24'd8955917, 24'd8697781, 24'd8378461, 24'd8061148, 24'd7808639, 24'd7670905, 24'd7675203, 24'd7820682, 24'd8078553, 24'd8397783, 24'd8715197, 24'd8967980, 24'd9106106, 24'd9102240, 24'd8957148, 24'd8699543, 24'd8380404, 24'd8062889, 24'd7809833, 24'd7671315, 24'd7674748, 24'd7819453, 24'd8076792, 24'd8395839, 24'd8713455, 24'd8966784, 24'd9105693, 24'd9102692, 24'd8958376, 24'd8701302, 
24'd8382348, 24'd8064632, 24'd7811030, 24'd7671730, 24'd7674298, 24'd7818227, 24'd8075034, 24'd8393896, 24'd8711711, 24'd8965585, 24'd9105276, 24'd9103140, 24'd8959599, 24'd8703060, 24'd8384291, 24'd8066377, 24'd7812231, 24'd7672150, 24'd7673854, 24'd7817006, 24'd8073277, 24'd8391952, 24'd8709965, 24'd8964381, 24'd9104854, 24'd9103582, 24'd8960818, 24'd8704815, 24'd8386235, 24'd8068124, 
24'd7813437, 24'd7672575, 24'd7673414, 24'd7815789, 24'd8071523, 24'd8390008, 24'd8708216, 24'd8963174, 24'd9104426, 24'd9104019, 24'd8962033, 24'd8706568, 24'd8388178, 24'd8069874, 24'd7814646, 24'd7673004, 24'd7672979, 24'd7814576, 24'd8069772, 24'd8388065, 24'd8706465, 24'd8961963, 24'd9103994, 24'd9104451, 24'd8963245, 24'd8708318, 24'd8390122, 24'd8071626, 24'd7815860, 24'd7673439, 
24'd7672550, 24'd7813366, 24'd8068022, 24'd8386121, 24'd8704712, 24'd8960747, 24'd9103556, 24'd9104878, 24'd8964452, 24'd8710067, 24'd8392065, 24'd8073380, 24'd7817077, 24'd7673879, 24'd7672125, 24'd7812161, 24'd8066275, 24'd8384178, 24'd8702957, 24'd8959527, 24'd9103114, 24'd9105300, 24'd8965655, 24'd8711813, 24'd8394009, 24'd8075136, 24'd7818299, 24'd7674324, 24'd7671705, 24'd7810960, 
24'd8064530, 24'd8382234, 24'd8701200, 24'd8958304, 24'd9102666, 24'd9105718, 24'd8966854, 24'd8713557, 24'd8395953, 24'd8076895, 24'd7819524, 24'd7674774, 24'd7671291, 24'd7809763, 24'd8062787, 24'd8380291, 24'd8699440, 24'd8957076, 24'd9102214, 24'd9106130, 24'd8968049, 24'd8715298, 24'd8397896, 24'd8078655, 24'd7820754, 24'd7675229, 24'd7670881, 24'd7808570, 24'd8061047, 24'd8378347, 
24'd8697678, 24'd8955845, 24'd9101756, 24'd9106537, 24'd8969240, 24'd8717038, 24'd8399839, 24'd8080418, 24'd7821987, 24'd7675689, 24'd7670477, 24'd7807381, 24'd8059309, 24'd8376404, 24'd8695914, 24'd8954609, 24'd9101294, 24'd9106939, 24'd8970427, 24'd8718775, 24'd8401783, 24'd8082183, 24'd7823225, 24'd7676154, 24'd7670077, 24'd7806196, 24'd8057573, 24'd8374461, 24'd8694148, 24'd8953370, 
24'd9100826, 24'd9107336, 24'd8971610, 24'd8720509, 24'd8403726, 24'd8083951, 24'd7824466, 24'd7676624, 24'd7669683, 24'd7805015, 24'd8055839, 24'd8372518, 24'd8692380, 24'd8952127, 24'd9100354, 24'd9107728, 24'd8972789, 24'd8722242, 24'd8405669, 24'd8085720, 24'd7825712, 24'd7677099, 24'd7669293, 24'd7803838, 24'd8054108, 24'd8370574, 24'd8690610, 24'd8950879, 24'd9099876, 24'd9108114, 
24'd8973964, 24'd8723972, 24'd8407612, 24'd8087491, 24'd7826961, 24'd7677579, 24'd7668909, 24'd7802666, 24'd8052379, 24'd8368632, 24'd8688837, 24'd8949628, 24'd9099394, 24'd9108496, 24'd8975134, 24'd8725699, 24'd8409555, 24'd8089265, 24'd7828214, 24'd7678064, 24'd7668530, 24'd7801497, 24'd8050653, 24'd8366689, 24'd8687063, 24'd8948373, 24'd9098906, 24'd9108873, 24'd8976301, 24'd8727425, 
24'd8411498, 24'd8091040, 24'd7829471, 24'd7678554, 24'd7668155, 24'd7800333, 24'd8048928, 24'd8364746, 24'd8685286, 24'd8947114, 24'd9098414, 24'd9109245, 24'd8977463, 24'd8729148, 24'd8413440, 24'd8092818, 24'd7830732, 24'd7679049, 24'd7667786, 24'd7799172, 24'd8047207, 24'd8362804, 24'd8683507, 24'd8945850, 24'd9097916, 24'd9109612, 24'd8978621, 24'd8730868, 24'd8415382, 24'd8094598, 
24'd7831998, 24'd7679549, 24'd7667422, 24'd7798016, 24'd8045487, 24'd8360861, 24'd8681726, 24'd8944584, 24'd9097414, 24'd9109973, 24'd8979775, 24'd8732586, 24'd8417325, 24'd8096380, 24'd7833266, 24'd7680054, 24'd7667063, 24'd7796864, 24'd8043770, 24'd8358919, 24'd8679943, 24'd8943313, 24'd9096907, 24'd9110330, 24'd8980925, 24'd8734302, 24'd8419267, 24'd8098164, 24'd7834539, 24'd7680564, 
24'd7666709, 24'd7795716, 24'd8042056, 24'd8356977, 24'd8678158, 24'd8942038, 24'd9096394, 24'd9110681, 24'd8982071, 24'd8736015, 24'd8421208, 24'd8099950, 24'd7835816, 24'd7681079, 24'd7666360, 24'd7794573, 24'd8040344, 24'd8355036, 24'd8676371, 24'd8940759, 24'd9095877, 24'd9111028, 24'd8983213, 24'd8737726, 24'd8423150, 24'd8101738, 24'd7837097, 24'd7681598, 24'd7666016, 24'd7793433, 
24'd8038634, 24'd8353094, 24'd8674582, 24'd8939477, 24'd9095355, 24'd9111369, 24'd8984350, 24'd8739435, 24'd8425091, 24'd8103528, 24'd7838381, 24'd7682123, 24'd7665677, 24'd7792298, 24'd8036927, 24'd8351153, 24'd8672791, 24'd8938190, 24'd9094828, 24'd9111705, 24'd8985483, 24'd8741141, 24'd8427032, 24'd8105320, 24'd7839669, 24'd7682653, 24'd7665343, 24'd7791167, 24'd8035222, 24'd8349212, 
24'd8670998, 24'd8936900, 24'd9094296, 24'd9112037, 24'd8986612, 24'd8742844, 24'd8428973, 24'd8107114, 24'd7840962, 24'd7683187, 24'd7665015, 24'd7790040, 24'd8033520, 24'd8347272, 24'd8669204, 24'd8935606, 24'd9093758, 24'd9112363, 24'd8987737, 24'd8744545, 24'd8430914, 24'd8108910, 24'd7842258, 24'd7683727, 24'd7664691, 24'd7788917, 24'd8031820, 24'd8345331, 24'd8667407, 24'd8934308, 
24'd9093216, 24'd9112684, 24'd8988858, 24'd8746244, 24'd8432854, 24'd8110708, 24'd7843557, 24'd7684271, 24'd7664372, 24'd7787798, 24'd8030123, 24'd8343391, 24'd8665608, 24'd8933006, 24'd9092669, 24'd9113000, 24'd8989975, 24'd8747940, 24'd8434794, 24'd8112507, 24'd7844861, 24'd7684821, 24'd7664059, 24'd7786684, 24'd8028428, 24'd8341451, 24'd8663807, 24'd8931701, 24'd9092118, 24'd9113311, 
24'd8991087, 24'd8749633, 24'd8436733, 24'd8114309, 24'd7846168, 24'd7685375, 24'd7663751, 24'd7785574, 24'd8026736, 24'd8339512, 24'd8662004, 24'd8930391, 24'd9091561, 24'd9113617, 24'd8992195, 24'd8751324, 24'd8438672, 24'd8116113, 24'd7847480, 24'd7685935, 24'd7663447, 24'd7784468, 24'd8025046, 24'd8337573, 24'd8660199, 24'd8929078, 24'd9090999, 24'd9113918, 24'd8993299, 24'd8753013, 
24'd8440611, 24'd8117919, 24'd7848795, 24'd7686499, 24'd7663149, 24'd7783366, 24'd8023359, 24'd8335634, 24'd8658393, 24'd8927761, 24'd9090432, 24'd9114213, 24'd8994398, 24'd8754698, 24'd8442550, 24'd8119726, 24'd7850114, 24'd7687068, 24'd7662856, 24'd7782269, 24'd8021675, 24'd8333696, 24'd8656584, 24'd8926441, 24'd9089861, 24'd9114504, 24'd8995494, 24'd8756382, 24'd8444488, 24'd8121536, 
24'd7851436, 24'd7687642, 24'd7662568, 24'd7781175, 24'd8019993, 24'd8331758, 24'd8654774, 24'd8925116, 24'd9089284, 24'd9114789, 24'd8996585, 24'd8758062, 24'd8446426, 24'd8123347, 24'd7852763, 24'd7688221, 24'd7662285, 24'd7780086, 24'd8018313, 24'd8329821, 24'd8652962, 24'd8923788, 24'd9088703, 24'd9115070, 24'd8997672, 24'd8759741, 24'd8448363, 24'd8125160, 24'd7854093, 24'd7688805, 
24'd7662007, 24'd7779002, 24'd8016636, 24'd8327883, 24'd8651148, 24'd8922456, 24'd9088116, 24'd9115345, 24'd8998754, 24'd8761416, 24'd8450300, 24'd8126975, 24'd7855427, 24'd7689394, 24'd7661734, 24'd7777921, 24'd8014962, 24'd8325947, 24'd8649332, 24'd8921120, 24'd9087525, 24'd9115615, 24'd8999832, 24'd8763089, 24'd8452236, 24'd8128792, 24'd7856764, 24'd7689988, 24'd7661466, 24'd7776845, 
24'd8013291, 24'd8324010, 24'd8647514, 24'd8919780, 24'd9086929, 24'd9115881, 24'd9000906, 24'd8764759, 24'd8454172, 24'd8130611, 24'd7858106, 24'd7690586, 24'd7661204, 24'd7775773, 24'd8011622, 24'd8322075, 24'd8645694, 24'd8918437, 24'd9086328, 24'd9116141, 24'd9001976, 24'd8766427, 24'd8456108, 24'd8132431, 24'd7859451, 24'd7691190, 24'd7660946, 24'd7774706, 24'd8009955, 24'd8320139, 
24'd8643873, 24'd8917090, 24'd9085722, 24'd9116396, 24'd9003041, 24'd8768092, 24'd8458043, 24'd8134253, 24'd7860800, 24'd7691798, 24'd7660694, 24'd7773643, 24'd8008292, 24'd8318204, 24'd8642050, 24'd8915740, 24'd9085111, 24'd9116645, 24'd9004102, 24'd8769754, 24'd8459978, 24'd8136077, 24'd7862152, 24'd7692411, 24'd7660447, 24'd7772584, 24'd8006631, 24'd8316270, 24'd8640225, 24'd8914385, 
24'd9084495, 24'd9116890, 24'd9005159, 24'd8771414, 24'd8461912, 24'd8137903, 24'd7863508, 24'd7693030, 24'd7660204, 24'd7771529, 24'd8004972, 24'd8314336, 24'd8638398, 24'd8913027, 24'd9083875, 24'd9117130, 24'd9006212, 24'd8773071, 24'd8463846, 24'd8139731, 24'd7864868, 24'd7693653, 24'd7659967, 24'd7770479, 24'd8003317, 24'd8312403, 24'd8636570, 24'd8911666, 24'd9083249, 24'd9117364, 
24'd9007260, 24'd8774725, 24'd8465779, 24'd8141560, 24'd7866232, 24'd7694280, 24'd7659735, 24'd7769433, 24'd8001664, 24'd8310470, 24'd8634740, 24'd8910300, 24'd9082619, 24'd9117594, 24'd9008304, 24'd8776377, 24'd8467711, 24'd8143391, 24'd7867599, 24'd7694913, 24'd7659509, 24'd7768391, 24'd8000013, 24'd8308538, 24'd8632908, 24'd8908931, 24'd9081984, 24'd9117818, 24'd9009343, 24'd8778026, 
24'd8469643, 24'd8145224, 24'd7868970, 24'd7695551, 24'd7659287, 24'd7767354, 24'd7998366, 24'd8306606, 24'd8631074, 24'd8907559, 24'd9081343, 24'd9118037, 24'd9010378, 24'd8779672, 24'd8471574, 24'd8147058, 24'd7870344, 24'd7696193, 24'd7659070, 24'd7766321, 24'd7996721, 24'd8304675, 24'd8629239, 24'd8906182, 24'd9080698, 24'd9118251, 24'd9011409, 24'd8781315, 24'd8473505, 24'd8148894, 
24'd7871722, 24'd7696841, 24'd7658859, 24'd7765293, 24'd7995079, 24'd8302744, 24'd8627402, 24'd8904802, 24'd9080049, 24'd9118460, 24'd9012435, 24'd8782956, 24'd8475436, 24'd8150732, 24'd7873104, 24'd7697493, 24'd7658652, 24'd7764268, 24'd7993440, 24'd8300815, 24'd8625563, 24'd8903419, 24'd9079394, 24'd9118664, 24'd9013457, 24'd8784594, 24'd8477365, 24'd8152572, 24'd7874489, 24'd7698150, 
24'd7658451, 24'd7763249, 24'd7991804, 24'd8298885, 24'd8623723, 24'd8902032, 24'd9078735, 24'd9118863, 24'd9014475, 24'd8786229, 24'd8479294, 24'd8154413, 24'd7875878, 24'd7698812, 24'd7658255, 24'd7762233, 24'd7990170, 24'd8296957, 24'd8621881, 24'd8900641, 24'd9078070, 24'd9119056, 24'd9015488, 24'd8787861, 24'd8481223, 24'd8156256, 24'd7877271, 24'd7699479, 24'd7658064, 24'd7761222, 
24'd7988539, 24'd8295029, 24'd8620037, 24'd8899246, 24'd9077401, 24'd9119245, 24'd9016497, 24'd8789490, 24'd8483150, 24'd8158100, 24'd7878667, 24'd7700150, 24'd7657878, 24'd7760216, 24'd7986911, 24'd8293101, 24'd8618192, 24'd8897848, 24'd9076727, 24'd9119428, 24'd9017501, 24'd8791117, 24'd8485077, 24'd8159946, 24'd7880067, 24'd7700827, 24'd7657697, 24'd7759213, 24'd7985286, 24'd8291174, 
24'd8616345, 24'd8896447, 24'd9076048, 24'd9119606, 24'd9018501, 24'd8792741, 24'd8487004, 24'd8161794, 24'd7881470, 24'd7701508, 24'd7657521, 24'd7758216, 24'd7983663, 24'd8289248, 24'd8614497, 24'd8895042, 24'd9075365, 24'd9119779, 24'd9019497, 24'd8794362, 24'd8488929, 24'd8163643, 24'd7882877, 24'd7702194, 24'd7657351, 24'd7757222, 24'd7982043, 24'd8287323, 24'd8612647, 24'd8893633, 
24'd9074676, 24'd9119947, 24'd9020488, 24'd8795980, 24'd8490854, 24'd8165494, 24'd7884287, 24'd7702885, 24'd7657185, 24'd7756233, 24'd7980427, 24'd8285398, 24'd8610795, 24'd8892221, 24'd9073983, 24'd9120110, 24'd9021475, 24'd8797596, 24'd8492779, 24'd8167346, 24'd7885701, 24'd7703580, 24'd7657025, 24'd7755249, 24'd7978813, 24'd8283474, 24'd8608942, 24'd8890805, 24'd9073285, 24'd9120268, 
24'd9022457, 24'd8799208, 24'd8494702, 24'd8169200, 24'd7887119, 24'd7704281, 24'd7656870, 24'd7754269, 24'd7977202, 24'd8281551, 24'd8607087, 24'd8889386, 24'd9072582, 24'd9120421, 24'd9023435, 24'd8800818, 24'd8496625, 24'd8171056, 24'd7888540, 24'd7704986, 24'd7656720, 24'd7753293, 24'd7975594, 24'd8279629, 24'd8605231, 24'd8887963, 24'd9071874, 24'd9120568, 24'd9024408, 24'd8802424, 
24'd8498547, 24'd8172913, 24'd7889964, 24'd7705696, 24'd7656575, 24'd7752322, 24'd7973988, 24'd8277707, 24'd8603373, 24'd8886537, 24'd9071162, 24'd9120710, 24'd9025377, 24'd8804028, 24'd8500468, 24'd8174771, 24'd7891392, 24'd7706411, 24'd7656435, 24'd7751355, 24'd7972386, 24'd8275786, 24'd8601514, 24'd8885108, 24'd9070445, 24'd9120848, 24'd9026342, 24'd8805629, 24'd8502389, 24'd8176631, 
24'd7892824, 24'd7707131, 24'd7656301, 24'd7750393, 24'd7970787, 24'd8273866, 24'd8599653, 24'd8883674, 24'd9069723, 24'd9120980, 24'd9027302, 24'd8807227, 24'd8504308, 24'd8178493, 24'd7894259, 24'd7707855, 24'd7656171, 24'd7749435, 24'd7969190, 24'd8271947, 24'd8597791, 24'd8882238, 24'd9068996, 24'd9121107, 24'd9028257, 24'd8808822, 24'd8506227, 24'd8180356, 24'd7895697, 24'd7708584, 
24'd7656047, 24'd7748482, 24'd7967597, 24'd8270029, 24'd8595927, 24'd8880798, 24'd9068264, 24'd9121228, 24'd9029208, 24'd8810414, 24'd8508145, 24'd8182220, 24'd7897139, 24'd7709318, 24'd7655928, 24'd7747533, 24'd7966006, 24'd8268111, 24'd8594062, 24'd8879354, 24'd9067528, 24'd9121345, 24'd9030155, 24'd8812003, 24'd8510063, 24'd8184086, 24'd7898584, 24'd7710057, 24'd7655814, 24'd7746589, 
24'd7964418, 24'd8266194, 24'd8592195, 24'd8877907, 24'd9066787, 24'd9121457, 24'd9031097, 24'd8813589, 24'd8511979, 24'd8185953, 24'd7900033, 24'd7710800, 24'd7655705, 24'd7745649, 24'd7962834, 24'd8264278, 24'd8590327, 24'd8876456, 24'd9066041, 24'd9121563, 24'd9032034, 24'd8815173, 24'd8513894, 24'd8187822, 24'd7901485, 24'd7711549, 24'd7655601, 24'd7744714, 24'd7961252, 24'd8262363, 
24'd8588458, 24'd8875003, 24'd9065291, 24'd9121664, 24'd9032967, 24'd8816753, 24'd8515809, 24'd8189692, 24'd7902941, 24'd7712302, 24'd7655502, 24'd7743783, 24'd7959673, 24'd8260449, 24'd8586587, 24'd8873545, 24'd9064535, 24'd9121760, 24'd9033896, 24'd8818330, 24'd8517723, 24'd8191564, 24'd7904400, 24'd7713059, 24'd7655409, 24'd7742857, 24'd7958098, 24'd8258536, 24'd8584715, 24'd8872085, 
24'd9063775, 24'd9121851, 24'd9034820, 24'd8819904, 24'd8519636, 24'd8193437, 24'd7905862, 24'd7713822, 24'd7655320, 24'd7741935, 24'd7956525, 24'd8256623, 24'd8582841, 24'd8870621, 24'd9063010, 24'd9121937, 24'd9035739, 24'd8821475, 24'd8521547, 24'd8195311, 24'd7907328, 24'd7714589, 24'd7655237, 24'd7741018, 24'd7954955, 24'd8254712, 24'd8580966, 24'd8869153, 24'd9062241, 24'd9122018, 
24'd9036654, 24'd8823043, 24'd8523458, 24'd8197187, 24'd7908797, 24'd7715361, 24'd7655159, 24'd7740105, 24'd7953389, 24'd8252801, 24'd8579090, 24'd8867682, 24'd9061467, 24'd9122093, 24'd9037565, 24'd8824608, 24'd8525368, 24'd8199064, 24'd7910269, 24'd7716137, 24'd7655086, 24'd7739197, 24'd7951825, 24'd8250892, 24'd8577212, 24'd8866208, 24'd9060688, 24'd9122164, 24'd9038470, 24'd8826170, 
24'd8527278, 24'd8200942, 24'd7911745, 24'd7716919, 24'd7655018, 24'd7738293, 24'd7950265, 24'd8248983, 24'd8575333, 24'd8864731, 24'd9059904, 24'd9122229, 24'd9039372, 24'd8827729, 24'd8529186, 24'd8202822, 24'd7913225, 24'd7717705, 24'd7654955, 24'd7737394, 24'd7948707, 24'd8247076, 24'd8573453, 24'd8863250, 24'd9059115, 24'd9122289, 24'd9040268, 24'd8829285, 24'd8531093, 24'd8204703, 
24'd7914707, 24'd7718495, 24'd7654898, 24'd7736500, 24'd7947153, 24'd8245169, 24'd8571571, 24'd8861765, 24'd9058322, 24'd9122344, 24'd9041161, 24'd8830838, 24'd8532999, 24'd8206585, 24'd7916193, 24'd7719291, 24'd7654845, 24'd7735610, 24'd7945602, 24'd8243264, 24'd8569689, 24'd8860278, 24'd9057525, 24'd9122394, 24'd9042048, 24'd8832388, 24'd8534904, 24'd8208468, 24'd7917682, 24'd7720091, 
24'd7654798, 24'd7734725, 24'd7944054, 24'd8241359, 24'd8567804, 24'd8858787, 24'd9056722, 24'd9122438, 24'd9042931, 24'd8833934, 24'd8536808, 24'd8210353, 24'd7919175, 24'd7720896, 24'd7654756, 24'd7733844, 24'd7942509, 24'd8239455, 24'd8565919, 24'd8857293, 24'd9055915, 24'd9122478, 24'd9043809, 24'd8835478, 24'd8538711, 24'd8212239, 24'd7920670, 24'd7721705, 24'd7654719, 24'd7732968, 
24'd7940967, 24'd8237553, 24'd8564032, 24'd8855796, 24'd9055103, 24'd9122512, 24'd9044683, 24'd8837018, 24'd8540613, 24'd8214126, 24'd7922169, 24'd7722520, 24'd7654687, 24'd7732097, 24'd7939428, 24'd8235651, 24'd8562144, 24'd8854295, 24'd9054287, 24'd9122542, 24'd9045552, 24'd8838555, 24'd8542514, 24'd8216015, 24'd7923672, 24'd7723338, 24'd7654661, 24'd7731230, 24'd7937893, 24'd8233751, 
24'd8560255, 24'd8852791, 24'd9053465, 24'd9122566, 24'd9046417, 24'd8840089, 24'd8544414, 24'd8217905, 24'd7925177, 24'd7724162, 24'd7654639, 24'd7730367, 24'd7936360, 24'd8231852, 24'd8558365, 24'd8851284, 24'd9052640, 24'd9122585, 24'd9047277, 24'd8841620, 24'd8546312, 24'd8219795, 24'd7926686, 24'd7724990, 24'd7654623, 24'd7729510, 24'd7934831, 24'd8229954, 24'd8556474, 24'd8849773, 
24'd9051809, 24'd9122598, 24'd9048132, 24'd8843148, 24'd8548210, 24'd8221688, 24'd7928198, 24'd7725823, 24'd7654612, 24'd7728657, 24'd7933305, 24'd8228057, 24'd8554581, 24'd8848260, 24'd9050974, 24'd9122607, 24'd9048983, 24'd8844672, 24'd8550107, 24'd8223581, 24'd7929713, 24'd7726660, 24'd7654605, 24'd7727808, 24'd7931782, 24'd8226161, 24'd8552687, 24'd8846743, 24'd9050134, 24'd9122611, 
24'd9049829, 24'd8846193, 24'd8552002, 24'd8225475, 24'd7931232, 24'd7727503, 24'd7654605, 24'd7726964, 24'd7930262, 24'd8224266, 24'd8550792, 24'd8845223, 24'd9049290, 24'd9122609, 24'd9050671, 24'd8847711, 24'd8553896, 24'd8227371, 24'd7932754, 24'd7728349, 24'd7654609, 24'd7726125, 24'd7928746, 24'd8222372, 24'd8548896, 24'd8843699, 24'd9048441, 24'd9122602, 24'd9051508, 24'd8849226, 
24'd8555789, 24'd8229267, 24'd7934279, 24'd7729201, 24'd7654618, 24'd7725291, 24'd7927233, 24'd8220480, 24'd8546999, 24'd8842173, 24'd9047587, 24'd9122590, 24'd9052340, 24'd8850738, 24'd8557681, 24'd8231165, 24'd7935807, 24'd7730057, 24'd7654633, 24'd7724461, 24'd7925723, 24'd8218588, 24'd8545101, 24'd8840643, 24'd9046729, 24'd9122573, 24'd9053167, 24'd8852246, 24'd8559572, 24'd8233064, 
24'd7937338, 24'd7730917, 24'd7654652, 24'd7723636, 24'd7924216, 24'd8216698, 24'd8543201, 24'd8839110, 24'd9045866, 24'd9122551, 24'd9053990, 24'd8853751, 24'd8561461, 24'd8234964, 24'd7938872, 24'd7731783, 24'd7654677, 24'd7722815, 24'd7922712, 24'd8214809, 24'd8541301, 24'd8837574, 24'd9044998, 24'd9122524, 24'd9054808, 24'd8855253, 24'd8563350, 24'd8236865, 24'd7940410, 24'd7732652, 
24'd7654707, 24'd7721999, 24'd7921212, 24'd8212922, 24'd8539399, 24'd8836035, 24'd9044126, 24'd9122491, 24'd9055622, 24'd8856752, 24'd8565237, 24'd8238767, 24'd7941951, 24'd7733527, 24'd7654742, 24'd7721188, 24'd7919715, 24'd8211035, 24'd8537496, 24'd8834493, 24'd9043249, 24'd9122453, 24'd9056431, 24'd8858247, 24'd8567123, 24'd8240670, 24'd7943495, 24'd7734406, 24'd7654782, 24'd7720382, 
24'd7918221, 24'd8209150, 24'd8535593, 24'd8832947, 24'd9042368, 24'd9122411, 24'd9057235, 24'd8859739, 24'd8569007, 24'd8242575, 24'd7945042, 24'd7735289, 24'd7654828, 24'd7719580, 24'd7916731, 24'd8207266, 24'd8533688, 24'd8831399, 24'd9041482, 24'd9122363, 24'd9058034, 24'd8861228, 24'd8570891, 24'd8244480, 24'd7946592, 24'd7736178, 24'd7654878, 24'd7718783, 24'd7915244, 24'd8205383, 
24'd8531782, 24'd8829847, 24'd9040592, 24'd9122310, 24'd9058829, 24'd8862713, 24'd8572773, 24'd8246386, 24'd7948145, 24'd7737070, 24'd7654934, 24'd7717990, 24'd7913760, 24'd8203502, 24'd8529875, 24'd8828292, 24'd9039696, 24'd9122251, 24'd9059619, 24'd8864195, 24'd8574653, 24'd8248293, 24'd7949701, 24'd7737968, 24'd7654995, 24'd7717202, 24'd7912280, 24'd8201622, 24'd8527968, 24'd8826735, 
24'd9038797, 24'd9122188, 24'd9060405, 24'd8865674, 24'd8576533, 24'd8250202, 24'd7951261, 24'd7738870, 24'd7655061, 24'd7716419, 24'd7910803, 24'd8199743, 24'd8526059, 24'd8825174, 24'd9037893, 24'd9122119, 24'd9061185, 24'd8867149, 24'd8578411, 24'd8252111, 24'd7952823, 24'd7739776, 24'd7655132, 24'd7715641, 24'd7909329, 24'd8197865, 24'd8524149, 24'd8823610, 24'd9036984, 24'd9122046, 
24'd9061961, 24'd8868622, 24'd8580288, 24'd8254021, 24'd7954388, 24'd7740687, 24'd7655208, 24'd7714867, 24'd7907859, 24'd8195989, 24'd8522239, 24'd8822043, 24'd9036071, 24'd9121967, 24'd9062733, 24'd8870090, 24'd8582163, 24'd8255932, 24'd7955957, 24'd7741603, 24'd7655289, 24'd7714099, 24'd7906392, 24'd8194115, 24'd8520327, 24'd8820473, 24'd9035153, 24'd9121883, 24'd9063499, 24'd8871555, 
24'd8584037, 24'd8257844, 24'd7957529, 24'd7742523, 24'd7655376, 24'd7713334, 24'd7904928, 24'd8192241, 24'd8518415, 24'd8818900, 24'd9034230, 24'd9121794, 24'd9064261, 24'd8873017, 24'd8585910, 24'd8259757, 24'd7959103, 24'd7743447, 24'd7655468, 24'd7712575, 24'd7903468, 24'd8190369, 24'd8516501, 24'd8817323, 24'd9033304, 24'd9121700, 24'd9065018, 24'd8874476, 24'd8587781, 24'd8261671, 
24'd7960681, 24'd7744377, 24'd7655564, 24'd7711820, 24'd7902011, 24'd8188498, 24'd8514587, 24'd8815744, 24'd9032372, 24'd9121600, 24'd9065770, 24'd8875931, 24'd8589651, 24'd8263586, 24'd7962261, 24'd7745310, 24'd7655666, 24'd7711070, 24'd7900558, 24'd8186629, 24'd8512672, 24'd8814162, 24'd9031436, 24'd9121496, 24'd9066518, 24'd8877383, 24'd8591520, 24'd8265501, 24'd7963845, 24'd7746248, 
24'd7655774, 24'd7710325, 24'd7899108, 24'd8184761, 24'd8510756, 24'd8812577, 24'd9030496, 24'd9121386, 24'd9067261, 24'd8878831, 24'd8593387, 24'd8267418, 24'd7965431, 24'd7747191, 24'd7655886, 24'd7709585, 24'd7897661, 24'd8182895, 24'd8508839, 24'd8810989, 24'd9029551, 24'd9121271, 24'd9067999, 24'd8880276, 24'd8595253, 24'd8269335, 24'd7967021, 24'd7748138, 24'd7656003, 24'd7708849, 
24'd7896218, 24'd8181030, 24'd8506921, 24'd8809398, 24'd9028602, 24'd9121151, 24'd9068732, 24'd8881717, 24'd8597117, 24'd8271253, 24'd7968613, 24'd7749090, 24'd7656126, 24'd7708118, 24'd7894778, 24'd8179166, 24'd8505003, 24'd8807804, 24'd9027648, 24'd9121026, 24'd9069460, 24'd8883155, 24'd8598980, 24'd8273172, 24'd7970209, 24'd7750046, 24'd7656253, 24'd7707392, 24'd7893342, 24'd8177304, 
24'd8503083, 24'd8806207, 24'd9026689, 24'd9120896, 24'd9070184, 24'd8884590, 24'd8600841, 24'd8275092, 24'd7971807, 24'd7751007, 24'd7656386, 24'd7706671, 24'd7891909, 24'd8175444, 24'd8501163, 24'd8804607, 24'd9025726, 24'd9120761, 24'd9070903, 24'd8886021, 24'd8602701, 24'd8277012, 24'd7973409, 24'd7751972, 24'd7656524, 24'd7705954, 24'd7890480, 24'd8173585, 24'd8499242, 24'd8803005, 
24'd9024759, 24'd9120620, 24'd9071617, 24'd8887448, 24'd8604559, 24'd8278934, 24'd7975013, 24'd7752941, 24'd7656667, 24'd7705242, 24'd7889055, 24'd8171727, 24'd8497320, 24'd8801399, 24'd9023787, 24'd9120475, 24'd9072327, 24'd8888872, 24'd8606416, 24'd8280856, 24'd7976620, 24'd7753915, 24'd7656815, 24'd7704535, 24'd7887632, 24'd8169871, 24'd8495398, 24'd8799791, 24'd9022811, 24'd9120324, 
24'd9073031, 24'd8890293, 24'd8608271, 24'd8282779, 24'd7978230, 24'd7754894, 24'd7656968, 24'd7703833, 24'd7886214, 24'd8168017, 24'd8493474, 24'd8798179, 24'd9021830, 24'd9120168, 24'd9073731, 24'd8891710, 24'd8610125, 24'd8284703, 24'd7979843, 24'd7755877, 24'd7657127, 24'd7703136, 24'd7884798, 24'd8166164, 24'd8491550, 24'd8796565, 24'd9020845, 24'd9120007, 24'd9074426, 24'd8893123, 
24'd8611977, 24'd8286627, 24'd7981458, 24'd7756864, 24'd7657290, 24'd7702443, 24'd7883387, 24'd8164312, 24'd8489626, 24'd8794948, 24'd9019856, 24'd9119841, 24'd9075116, 24'd8894533, 24'd8613828, 24'd8288552, 24'd7983077, 24'd7757856, 24'd7657459, 24'd7701755, 24'd7881979, 24'd8162463, 24'd8487700, 24'd8793328, 24'd9018862, 24'd9119670, 24'd9075802, 24'd8895939, 24'd8615677, 24'd8290478, 
24'd7984698, 24'd7758852, 24'd7657633, 24'd7701072, 24'd7880574, 24'd8160614, 24'd8485774, 24'd8791705, 24'd9017863, 24'd9119493, 24'd9076482, 24'd8897342, 24'd8617524, 24'd8292404, 24'd7986323, 24'd7759853, 24'd7657812, 24'd7700394, 24'd7879173, 24'd8158768, 24'd8483847, 24'd8790079, 24'd9016860, 24'd9119312, 24'd9077158, 24'd8898741, 24'd8619370, 24'd8294331, 24'd7987950, 24'd7760858, 
24'd7657996, 24'd7699721, 24'd7877775, 24'd8156923, 24'd8481920, 24'd8788451, 24'd9015853, 24'd9119125, 24'd9077829, 24'd8900137, 24'd8621214, 24'd8296259, 24'd7989580, 24'd7761867, 24'd7658185, 24'd7699053, 24'd7876382, 24'd8155079, 24'd8479992, 24'd8786819, 24'd9014842, 24'd9118933, 24'd9078495, 24'd8901529, 24'd8623057, 24'd8298188, 24'd7991212, 24'd7762881, 24'd7658379, 24'd7698389, 
24'd7874991, 24'd8153237, 24'd8478063, 24'd8785185, 24'd9013826, 24'd9118736, 24'd9079156, 24'd8902917, 24'd8624898, 24'd8300117, 24'd7992848, 24'd7763899, 24'd7658579, 24'd7697730, 24'd7873605, 24'd8151397, 24'd8476133, 24'd8783548, 24'd9012805, 24'd9118534, 24'd9079813, 24'd8904302, 24'd8626737, 24'd8302046, 24'd7994486, 24'd7764922, 24'd7658783, 24'd7697076, 24'd7872222, 24'd8149559, 
24'd8474203, 24'd8781909, 24'd9011780, 24'd9118327, 24'd9080464, 24'd8905684, 24'd8628575, 24'd8303977, 24'd7996127, 24'd7765949, 24'd7658993, 24'd7696427, 24'd7870842, 24'd8147722, 24'd8472273, 24'd8780266, 24'd9010751, 24'd9118115, 24'd9081111, 24'd8907061, 24'd8630411, 24'd8305908, 24'd7997771, 24'd7766980, 24'd7659208, 24'd7695783, 24'd7869466, 24'd8145887, 24'd8470342, 24'd8778621, 
24'd9009718, 24'd9117898, 24'd9081753, 24'd8908435, 24'd8632245, 24'd8307839, 24'd7999417, 24'd7768016, 24'd7659428, 24'd7695143, 24'd7868094, 24'd8144054, 24'd8468410, 24'd8776973, 24'd9008680, 24'd9117675, 24'd9082390, 24'd8909806, 24'd8634077, 24'd8309771, 24'd8001067, 24'd7769056, 24'd7659653, 24'd7694509, 24'd7866726, 24'd8142222, 24'd8466478, 24'd8775323, 24'd9007638, 24'd9117448, 
24'd9083022, 24'd8911172, 24'd8635908, 24'd8311704, 24'd8002719, 24'd7770100, 24'd7659883, 24'd7693879, 24'd7865361, 24'd8140392, 24'd8464545, 24'd8773669, 24'd9006591, 24'd9117215, 24'd9083649, 24'd8912535, 24'd8637737, 24'd8313637, 24'd8004373, 24'd7771149, 24'd7660118, 24'd7693254, 24'd7864000, 24'd8138564, 24'd8462611, 24'd8772013, 24'd9005540, 24'd9116977, 24'd9084271, 24'd8913895, 
24'd8639565, 24'd8315571, 24'd8006031, 24'd7772202, 24'd7660358, 24'd7692634, 24'd7862642, 24'd8136737, 24'd8460677, 24'd8770355, 24'd9004485, 24'd9116734, 24'd9084889, 24'd8915250, 24'd8641390, 24'd8317505, 24'd8007691, 24'd7773259, 24'd7660604, 24'd7692019, 24'd7861288, 24'd8134913, 24'd8458743, 24'd8768693, 24'd9003426, 24'd9116486, 24'd9085501, 24'd8916602, 24'd8643214, 24'd8319440, 
24'd8009353, 24'd7774321, 24'd7660854, 24'd7691409, 24'd7859938, 24'd8133090, 24'd8456808, 24'd8767029, 24'd9002362, 24'd9116233, 24'd9086109, 24'd8917951, 24'd8645036, 24'd8321375, 24'd8011019, 24'd7775387, 24'd7661110, 24'd7690804, 24'd7858592, 24'd8131269, 24'd8454873, 24'd8765363, 24'd9001294, 24'd9115975, 24'd9086712, 24'd8919295, 24'd8646856, 24'd8323310, 24'd8012687, 24'd7776457, 
24'd7661371, 24'd7690203, 24'd7857249, 24'd8129449, 24'd8452937, 24'd8763693, 24'd9000221, 24'd9115712, 24'd9087310, 24'd8920636, 24'd8648675, 24'd8325246, 24'd8014357, 24'd7777532, 24'd7661637, 24'd7689608, 24'd7855910, 24'd8127632, 24'd8451000, 24'd8762021, 24'd8999145, 24'd9115443, 24'd9087903, 24'd8921973, 24'd8650491, 24'd8327183, 24'd8016031, 24'd7778610, 24'd7661908, 24'd7689017, 
24'd7854575, 24'd8125816, 24'd8449064, 24'd8760347, 24'd8998064, 24'd9115170, 24'd9088491, 24'd8923306, 24'd8652306, 24'd8329120, 24'd8017706, 24'd7779694, 24'd7662184, 24'd7688432, 24'd7853243, 24'd8124002, 24'd8447126, 24'd8758670, 24'd8996978, 24'd9114891, 24'd9089074, 24'd8924636, 24'd8654119, 24'd8331057, 24'd8019385, 24'd7780781, 24'd7662465, 24'd7687851, 24'd7851916, 24'd8122190, 
24'd8445189, 24'd8756990, 24'd8995889, 24'd9114608, 24'd9089653, 24'd8925962, 24'd8655930, 24'd8332995, 24'd8021066, 24'd7781873, 24'd7662751, 24'd7687275, 24'd7850592, 24'd8120380, 24'd8443251, 24'd8755308, 24'd8994795, 24'd9114319, 24'd9090226, 24'd8927284, 24'd8657739, 24'd8334933, 24'd8022750, 24'd7782969, 24'd7663042, 24'd7686704, 24'd7849271, 24'd8118572, 24'd8441312, 24'd8753623, 
24'd8993697, 24'd9114025, 24'd9090794, 24'd8928602, 24'd8659546, 24'd8336872, 24'd8024436, 24'd7784069, 24'd7663339, 24'd7686138, 24'd7847955, 24'd8116766, 24'd8439374, 24'd8751935, 24'd8992595, 24'd9113726, 24'd9091358, 24'd8929917, 24'd8661352, 24'd8338811, 24'd8026125, 24'd7785173, 24'd7663640, 24'd7685577, 24'd7846642, 24'd8114961, 24'd8437435, 24'd8750245, 24'd8991488, 24'd9113422, 
24'd9091917, 24'd8931228, 24'd8663155, 24'd8340750, 24'd8027816, 24'd7786282, 24'd7663947, 24'd7685021, 24'd7845333, 24'd8113159, 24'd8435495, 24'd8748552, 24'd8990377, 24'd9113113, 24'd9092470, 24'd8932535, 24'd8664957, 24'd8342690, 24'd8029510, 24'd7787395, 24'd7664258, 24'd7684470, 24'd7844028, 24'd8111358, 24'd8433555, 24'd8746857, 24'd8989262, 24'd9112799, 24'd9093019, 24'd8933838, 
24'd8666756, 24'd8344630, 24'd8031206, 24'd7788512, 24'd7664575, 24'd7683923, 24'd7842727, 24'd8109560, 24'd8431615, 24'd8745160, 24'd8988143, 24'd9112480, 24'd9093563, 24'd8935137, 24'd8668554, 24'd8346570, 24'd8032905, 24'd7789633, 24'd7664897, 24'd7683382, 24'd7841430, 24'd8107763, 24'd8429675, 24'd8743460, 24'd8987020, 24'd9112155, 24'd9094102, 24'd8936432, 24'd8670350, 24'd8348510, 
24'd8034606, 24'd7790758, 24'd7665224, 24'd7682846, 24'd7840136, 24'd8105968, 24'd8427734, 24'd8741757, 24'd8985892, 24'd9111826, 24'd9094636, 24'd8937724, 24'd8672143, 24'd8350451, 24'd8036310, 24'd7791888, 24'd7665556, 24'd7682314, 24'd7838847, 24'd8104176, 24'd8425793, 24'd8740052, 24'd8984760, 24'd9111491, 24'd9095165, 24'd8939012, 24'd8673935, 24'd8352392, 24'd8038016, 24'd7793022, 
24'd7665893, 24'd7681788, 24'd7837561, 24'd8102385, 24'd8423852, 24'd8738344, 24'd8983624, 24'd9111152, 24'd9095689, 24'd8940296, 24'd8675725, 24'd8354334, 24'd8039725, 24'd7794160, 24'd7666235, 24'd7681266, 24'd7836279, 24'd8100596, 24'd8421911, 24'd8736634, 24'd8982484, 24'd9110807, 24'd9096208, 24'd8941576, 24'd8677512, 24'd8356275, 24'd8041436, 24'd7795302, 24'd7666582, 24'd7680749, 
24'd7835001, 24'd8098810, 24'd8419969, 24'd8734922, 24'd8981340, 24'd9110457, 24'd9096722, 24'd8942852, 24'd8679298, 24'd8358217, 24'd8043150, 24'd7796449, 24'd7666934, 24'd7680238, 24'd7833726, 24'd8097025, 24'd8418027, 24'd8733207, 24'd8980192, 24'd9110103, 24'd9097231, 24'd8944124, 24'd8681082, 24'd8360159, 24'd8044866, 24'd7797599, 24'd7667292, 24'd7679731, 24'd7832456, 24'd8095242, 
24'd8416085, 24'd8731490, 24'd8979039, 24'd9109743, 24'd9097735, 24'd8945393, 24'd8682863, 24'd8362101, 24'd8046585, 24'd7798754, 24'd7667654, 24'd7679229, 24'd7831190, 24'd8093462, 24'd8414143, 24'd8729770, 24'd8977882, 24'd9109378, 24'd9098235, 24'd8946657, 24'd8684643, 24'd8364044, 24'd8048306, 24'd7799913, 24'd7668021, 24'd7678733, 24'd7829927, 24'd8091683, 24'd8412200, 24'd8728048, 
24'd8976721, 24'd9109008, 24'd9098729, 24'd8947918, 24'd8686420, 24'd8365986, 24'd8050029, 24'd7801076, 24'd7668394, 24'd7678241, 24'd7828668, 24'd8089907, 24'd8410257, 24'd8726324, 24'd8975556, 24'd9108633, 24'd9099218, 24'd8949174, 24'd8688196, 24'd8367929, 24'd8051754, 24'd7802243, 24'd7668771, 24'd7677754, 24'd7827414, 24'd8088132, 24'd8408315, 24'd8724597, 24'd8974387, 24'd9108253, 
24'd9099702, 24'd8950427, 24'd8689969, 24'd8369872, 24'd8053482, 24'd7803414, 24'd7669154, 24'd7677272, 24'd7826163, 24'd8086360, 24'd8406372, 24'd8722868, 24'd8973214, 24'd9107868, 24'd9100182, 24'd8951676, 24'd8691740, 24'd8371815, 24'd8055213, 24'd7804589, 24'd7669541, 24'd7676796, 24'd7824916, 24'd8084590, 24'd8404429, 24'd8721136, 24'd8972037, 24'd9107478, 24'd9100656, 24'd8952921, 
24'd8693509, 24'd8373758, 24'd8056945, 24'd7805768, 24'd7669934, 24'd7676324, 24'd7823673, 24'd8082822, 24'd8402485, 24'd8719402, 24'd8970855, 24'd9107083, 24'd9101125, 24'd8954162, 24'd8695276, 24'd8375701, 24'd8058680, 24'd7806952, 24'd7670332, 24'd7675857, 24'd7822434, 24'd8081056, 24'd8400542, 24'd8717666, 24'd8969670, 24'd9106683, 24'd9101590, 24'd8955399, 24'd8697041, 24'd8377644, 
24'd8060418, 24'd7808139, 24'd7670734, 24'd7675395, 24'd7821199, 24'd8079293, 24'd8398599, 24'd8715928, 24'd8968480, 24'd9106277, 24'd9102049, 24'd8956632, 24'd8698803, 24'd8379588, 24'd8062157, 24'd7809331, 24'd7671142, 24'd7674938, 24'd7819968, 24'd8077531, 24'd8396655, 24'd8714187, 24'd8967287, 24'd9105867, 24'd9102503, 24'd8957860, 24'd8700564, 24'd8381531, 24'd8063899, 24'd7810526, 
24'd7671555, 24'd7674487, 24'd7818742, 24'd8075772, 24'd8394712, 24'd8712444, 24'd8966089, 24'd9105452, 24'd9102952, 24'd8959085, 24'd8702322, 24'd8383475, 24'd8065644, 24'd7811726, 24'd7671973, 24'd7674040, 24'd7817519, 24'd8074015, 24'd8392768, 24'd8710699, 24'd8964887, 24'd9105032, 24'd9103397, 24'd8960306, 24'd8704078, 24'd8385418, 24'd8067390, 24'd7812930, 24'd7672395, 24'd7673598, 
24'd7816300, 24'd8072260, 24'd8390825, 24'd8708951, 24'd8963682, 24'd9104606, 24'd9103836, 24'd8961523, 24'd8705832, 24'd8387362, 24'd8069139, 24'd7814138, 24'd7672823, 24'd7673161, 24'd7815085, 24'd8070507, 24'd8388881, 24'd8707201, 24'd8962472, 24'd9104176, 24'd9104270, 24'd8962736, 24'd8707583, 24'd8389306, 24'd8070890, 24'd7815350, 24'd7673256, 24'd7672729, 24'd7813874, 24'd8068757, 
24'd8386938, 24'd8705449, 24'd8961258, 24'd9103741, 24'd9104700, 24'd8963945, 24'd8709333, 24'd8391249, 24'd8072643, 24'd7816565, 24'd7673694, 24'd7672303, 24'd7812667, 24'd8067009, 24'd8384994, 24'd8703695, 24'd8960040, 24'd9103300, 24'd9105124, 24'd8965150, 24'd8711080, 24'd8393193, 24'd8074398, 24'd7817785, 24'd7674137, 24'd7671881, 24'd7811464, 24'd8065263, 24'd8383051, 24'd8701938, 
24'd8958818, 24'd9102855, 24'd9105543, 24'd8966351, 24'd8712825, 24'd8395136, 24'd8076156, 24'd7819009, 24'd7674585, 24'd7671464, 24'd7810265, 24'd8063519, 24'd8381107, 24'd8700180, 24'd8957593, 24'd9102404, 24'd9105957, 24'd8967548, 24'd8714567, 24'd8397080, 24'd8077916, 24'd7820237, 24'd7675038, 24'd7671053, 24'd7809070, 24'd8061777, 24'd8379164, 24'd8698419, 24'd8956363, 24'd9101949, 
24'd9106366, 24'd8968740, 24'd8716307, 24'd8399023, 24'd8079678, 24'd7821469, 24'd7675496, 24'd7670646, 24'd7807880, 24'd8060038, 24'd8377220, 24'd8696656, 24'd8955129, 24'd9101489, 24'd9106770, 24'd8969929, 24'd8718045, 24'd8400966, 24'd8081442, 24'd7822704, 24'd7675958, 24'd7670244, 24'd7806693, 24'd8058302, 24'd8375277, 24'd8694890, 24'd8953891, 24'd9101023, 24'd9107170, 24'd8971114, 
24'd8719781, 24'd8402910, 24'd8083208, 24'd7823944, 24'd7676426, 24'd7669848, 24'd7805511, 24'd8056567, 24'd8373334, 24'd8693123, 24'd8952649, 24'd9100553, 24'd9107564, 24'd8972294, 24'd8721514, 24'd8404853, 24'd8084976, 24'd7825188, 24'd7676899, 24'd7669456, 24'd7804332, 24'd8054835, 24'd8371391, 24'd8691354, 24'd8951404, 24'd9100077, 24'd9107953, 24'd8973471, 24'd8723245, 24'd8406796, 
24'd8086747, 24'd7826436, 24'd7677377, 24'd7669070, 24'd7803158, 24'd8053105, 24'd8369448, 24'd8689582, 24'd8950154, 24'd9099597, 24'd9108337, 24'd8974643, 24'd8724974, 24'd8408739, 24'd8088520, 24'd7827687, 24'd7677860, 24'd7668688, 24'd7801987, 24'd8051378, 24'd8367505, 24'd8687808, 24'd8948900, 24'd9099112, 24'd9108715, 24'd8975811, 24'd8726700, 24'd8410682, 24'd8090294, 24'd7828943, 
24'd7678348, 24'd7668312, 24'd7800821, 24'd8049652, 24'd8365562, 24'd8686032, 24'd8947643, 24'd9098621, 24'd9109089, 24'd8976975, 24'd8728424, 24'd8412624, 24'd8092071, 24'd7830202, 24'd7678841, 24'd7667941, 24'd7799659, 24'd8047930, 24'd8363620, 24'd8684255, 24'd8946382, 24'd9098126, 24'd9109458, 24'd8978135, 24'd8730146, 24'd8414567, 24'd8093850, 24'd7831466, 24'd7679339, 24'd7667574, 
24'd7798501, 24'd8046209, 24'd8361677, 24'd8682475, 24'd8945116, 24'd9097626, 24'd9109822, 24'd8979291, 24'd8731865, 24'd8416509, 24'd8095631, 24'd7832733, 24'd7679841, 24'd7667213, 24'd7797348, 24'd8044491, 24'd8359735, 24'd8680693, 24'd8943847, 24'd9097120, 24'd9110181, 24'd8980443, 24'd8733582, 24'd8418451, 24'd8097414, 24'd7834004, 24'd7680349, 24'd7666857, 24'd7796198, 24'd8042776, 
24'd8357793, 24'd8678908, 24'd8942574, 24'd9096610, 24'd9110534, 24'd8981590, 24'd8735296, 24'd8420393, 24'd8099199, 24'd7835279, 24'd7680862, 24'd7666506, 24'd7795053, 24'd8041063, 24'd8355851, 24'd8677122, 24'd8941297, 24'd9096095, 24'd9110883, 24'd8982734, 24'd8737008, 24'd8422334, 24'd8100986, 24'd7836558, 24'd7681379, 24'd7666160, 24'd7793911, 24'd8039352, 24'd8353910, 24'd8675334, 
24'd8940016, 24'd9095575, 24'd9111226, 24'd8983873, 24'd8738717, 24'd8424276, 24'd8102776, 24'd7837841, 24'd7681902, 24'd7665819, 24'd7792774, 24'd8037644, 24'd8351969, 24'd8673544, 24'd8938731, 24'd9095050, 24'd9111565, 24'd8985008, 24'd8740424, 24'd8426217, 24'd8104567, 24'd7839128, 24'd7682430, 24'd7665483, 24'd7791641, 24'd8035938, 24'd8350027, 24'd8671752, 24'd8937442, 24'd9094520, 
24'd9111898, 24'd8986139, 24'd8742129, 24'd8428158, 24'd8106360, 24'd7840418, 24'd7682962, 24'd7665152, 24'd7790512, 24'd8034235, 24'd8348087, 24'd8669958, 24'd8936150, 24'd9093985, 24'd9112226, 24'd8987265, 24'd8743831, 24'd8430099, 24'd8108155, 24'd7841713, 24'd7683500, 24'd7664826, 24'd7789388, 24'd8032534, 24'd8346146, 24'd8668162, 24'd8934854, 24'd9093445, 24'd9112550, 24'd8988388, 
24'd8745531, 24'd8432039, 24'd8109952, 24'd7843011, 24'd7684042, 24'd7664506, 24'd7788268, 24'd8030836, 24'd8344206, 24'd8666364, 24'd8933554, 24'd9092900, 24'd9112868, 24'd8989506, 24'd8747228, 24'd8433979, 24'd8111751, 24'd7844313, 24'd7684590, 24'd7664190, 24'd7787151, 24'd8029140, 24'd8342266, 24'd8664564, 24'd8932250, 24'd9092350, 24'd9113181, 24'd8990620, 24'd8748922, 24'd8435919, 
24'd8113552, 24'd7845619, 24'd7685142, 24'd7663879, 24'd7786039, 24'd8027447, 24'd8340327, 24'd8662762, 24'd8930942, 24'd9091795, 24'd9113489, 24'd8991730, 24'd8750614, 24'd8437858, 24'd8115355, 24'd7846928, 24'd7685699, 24'd7663574, 24'd7784932, 24'd8025756, 24'd8338388, 24'd8660958, 24'd8929630, 24'd9091235, 24'd9113792, 24'd8992836, 24'd8752304, 24'd8439797, 24'd8117160, 24'd7848242, 
24'd7686261, 24'd7663274, 24'd7783828, 24'd8024068, 24'd8336449, 24'd8659152, 24'd8928315, 24'd9090671, 24'd9114090, 24'd8993937, 24'd8753991, 24'd8441736, 24'd8118967, 24'd7849559, 24'd7686828, 24'd7662978, 24'd7782729, 24'd8022382, 24'd8334510, 24'd8657344, 24'd8926996, 24'd9090101, 24'd9114382, 24'd8995034, 24'd8755675, 24'd8443674, 24'd8120775, 24'd7850880, 24'd7687400, 24'd7662688, 
24'd7781634, 24'd8020699, 24'd8332572, 24'd8655535, 24'd8925673, 24'd9089527, 24'd9114670, 24'd8996127, 24'd8757357, 24'd8445612, 24'd8122586, 24'd7852205, 24'd7687977, 24'd7662403, 24'd7780543, 24'd8019018, 24'd8330634, 24'd8653723, 24'd8924346, 24'd9088947, 24'd9114953, 24'd8997216, 24'd8759036, 24'd8447549, 24'd8124398, 24'd7853534, 24'd7688559, 24'd7662123, 24'd7779457, 24'd8017340, 
24'd8328697, 24'd8651910, 24'd8923016, 24'd9088363, 24'd9115230, 24'd8998300, 24'd8760713, 24'd8449486, 24'd8126212, 24'd7854866, 24'd7689146, 24'd7661848, 24'd7778375, 24'd8015665, 24'd8326760, 24'd8650095, 24'd8921682, 24'd9087774, 24'd9115502, 24'd8999380, 24'd8762387, 24'd8451423, 24'd8128028, 24'd7856202, 24'd7689738, 24'd7661578, 24'd7777297, 24'd8013992, 24'd8324824, 24'd8648278, 
24'd8920344, 24'd9087180, 24'd9115770, 24'd9000456, 24'd8764058, 24'd8453359, 24'd8129846, 24'd7857542, 24'd7690334, 24'd7661313, 24'd7776223, 24'd8012322, 24'd8322888, 24'd8646459, 24'd8919002, 24'd9086581, 24'd9116032, 24'd9001527, 24'd8765727, 24'd8455295, 24'd8131666, 24'd7858885, 24'd7690936, 24'd7661054, 24'd7775154, 24'd8010655, 24'd8320952, 24'd8644638, 24'd8917657, 24'd9085977, 
24'd9116289, 24'd9002594, 24'd8767393, 24'd8457230, 24'd8133488, 24'd7860233, 24'd7691542, 24'd7660799, 24'd7774089, 24'd8008990, 24'd8319017, 24'd8642816, 24'd8916307, 24'd9085368, 24'd9116541, 24'd9003657, 24'd8769056, 24'd8459165, 24'd8135311, 24'd7861583, 24'd7692153, 24'd7660550, 24'd7773028, 24'd8007328, 24'd8317083, 24'd8640992, 24'd8914955, 24'd9084754, 24'd9116788, 24'd9004716, 
24'd8770717, 24'd8461100, 24'd8137136, 24'd7862938, 24'd7692769, 24'd7660306, 24'd7771971, 24'd8005669, 24'd8315148, 24'd8639166, 24'd8913598, 24'd9084136, 24'd9117030, 24'd9005770, 24'd8772375, 24'd8463033, 24'd8138963, 24'd7864296, 24'd7693390, 24'd7660066, 24'd7770919, 24'd8004012, 24'd8313215, 24'd8637338, 24'd8912238, 24'd9083512, 24'd9117266, 24'd9006820, 24'd8774031, 24'd8464967, 
24'd8140791, 24'd7865658, 24'd7694016, 24'd7659832, 24'd7769872, 24'd8002358, 24'd8311282, 24'd8635509, 24'd8910874, 24'd9082884, 24'd9117498, 24'd9007866, 24'd8775683, 24'd8466899, 24'd8142622, 24'd7867024, 24'd7694647, 24'd7659603, 24'd7768828, 24'd8000706, 24'd8309349, 24'd8633678, 24'd8909507, 24'd9082251, 24'd9117724, 24'd9008907, 24'd8777333, 24'd8468832, 24'd8144454, 24'd7868393, 
24'd7695282, 24'd7659379, 24'd7767789, 24'd7999058, 24'd8307417, 24'd8631845, 24'd8908136, 24'd9081613, 24'd9117946, 24'd9009944, 24'd8778981, 24'd8470763, 24'd8146287, 24'd7869766, 24'd7695923, 24'd7659161, 24'd7766754, 24'd7997412, 24'd8305486, 24'd8630010, 24'd8906761, 24'd9080970, 24'd9118162, 24'd9010976, 24'd8780625, 24'd8472694, 24'd8148123, 24'd7871143, 24'd7696568, 24'd7658947, 
24'd7765724, 24'd7995769, 24'd8303555, 24'd8628174, 24'd8905382, 24'd9080322, 24'd9118373, 24'd9012005, 24'd8782267, 24'd8474625, 24'd8149960, 24'd7872523, 24'd7697218, 24'd7658738, 24'd7764698, 24'd7994128, 24'd8301625, 24'd8626336, 24'd8904000, 24'd9079670, 24'd9118579, 24'd9013028, 24'd8783906, 24'd8476555, 24'd8151799, 24'd7873907, 24'd7697873, 24'd7658535, 24'd7763676, 24'd7992491, 
24'd8299696, 24'd8624496, 24'd8902615, 24'd9079012, 24'd9118780, 24'd9014048, 24'd8785542, 24'd8478484, 24'd8153639, 24'd7875295, 24'd7698533, 24'd7658337, 24'd7762659, 24'd7990856, 24'd8297767, 24'd8622655, 24'd8901225, 24'd9078350, 24'd9118976, 24'd9015063, 24'd8787176, 24'd8480413, 24'd8155481, 24'd7876686, 24'd7699198, 24'd7658143, 24'd7761646, 24'd7989224, 24'd8295838, 24'd8620812, 
24'd8899833, 24'd9077683, 24'd9119166, 24'd9016073, 24'd8788806, 24'd8482341, 24'd8157325, 24'd7878080, 24'd7699868, 24'd7657955, 24'd7760638, 24'd7987594, 24'd8293911, 24'd8618967, 24'd8898436, 24'd9077011, 24'd9119352, 24'd9017080, 24'd8790434, 24'd8484268, 24'd8159171, 24'd7879478, 24'd7700542, 24'd7657772, 24'd7759634, 24'd7985968, 24'd8291984, 24'd8617121, 24'd8897036, 24'd9076334, 
24'd9119532, 24'd9018082, 24'd8792059, 24'd8486195, 24'd8161018, 24'd7880880, 24'd7701221, 24'd7657595, 24'd7758634, 24'd7984344, 24'd8290057, 24'd8615273, 24'd8895633, 24'd9075652, 24'd9119707, 24'd9019079, 24'd8793682, 24'd8488121, 24'd8162866, 24'd7882286, 24'd7701905, 24'd7657422, 24'd7757639, 24'd7982723, 24'd8288132, 24'd8613424, 24'd8894225, 24'd9074966, 24'd9119878, 24'd9020072, 
24'd8795301, 24'd8490046, 24'd8164716, 24'd7883695, 24'd7702594, 24'd7657254, 24'd7756648, 24'd7981105, 24'd8286207, 24'd8611573, 24'd8892815, 24'd9074275, 24'd9120043, 24'd9021061, 24'd8796917, 24'd8491970, 24'd8166568, 24'd7885107, 24'd7703288, 24'd7657092, 24'd7755662, 24'd7979490, 24'd8284283, 24'd8609720, 24'd8891401, 24'd9073579, 24'd9120202, 24'd9022045, 24'd8798531, 24'd8493894, 
24'd8168421, 24'd7886523, 24'd7703986, 24'd7656935, 24'd7754680, 24'd7977878, 24'd8282359, 24'd8607866, 24'd8889983, 24'd9072878, 24'd9120357, 24'd9023025, 24'd8800142, 24'd8495817, 24'd8170276, 24'd7887942, 24'd7704689, 24'd7656782, 24'd7753702, 24'd7976269, 24'd8280436, 24'd8606011, 24'd8888562, 24'd9072172, 24'd9120507, 24'd9024000, 24'd8801750, 24'd8497740, 24'd8172133, 24'd7889365, 
24'd7705397, 24'd7656635, 24'd7752729, 24'd7974662, 24'd8278514, 24'd8604154, 24'd8887137, 24'd9071462, 24'd9120651, 24'd9024971, 24'd8803355, 24'd8499661, 24'd8173990, 24'd7890792, 24'd7706110, 24'd7656493, 24'd7751761, 24'd7973059, 24'd8276593, 24'd8602295, 24'd8885708, 24'd9070747, 24'd9120791, 24'd9025937, 24'd8804957, 24'd8501582, 24'd8175850, 24'd7892222, 24'd7706828, 24'd7656357, 
24'd7750797, 24'd7971458, 24'd8274673, 24'd8600435, 24'd8884277, 24'd9070027, 24'd9120925, 24'd9026899, 24'd8806556, 24'd8503502, 24'd8177711, 24'd7893655, 24'd7707550, 24'd7656225, 24'd7749837, 24'd7969860, 24'd8272753, 24'd8598573, 24'd8882842, 24'd9069302, 24'd9121054, 24'd9027856, 24'd8808152, 24'd8505421, 24'd8179573, 24'd7895092, 24'd7708277, 24'd7656098, 24'd7748882, 24'd7968266, 
24'd8270834, 24'd8596710, 24'd8881403, 24'd9068572, 24'd9121178, 24'd9028809, 24'd8809746, 24'd8507340, 24'd8181437, 24'd7896533, 24'd7709009, 24'd7655977, 24'd7747931, 24'd7966674, 24'd8268916, 24'd8594846, 24'd8879961, 24'd9067838, 24'd9121297, 24'd9029758, 24'd8811336, 24'd8509257, 24'd8183302, 24'd7897977, 24'd7709746, 24'd7655861, 24'd7746985, 24'd7965085, 24'd8266999, 24'd8592980, 
24'd8878515, 24'd9067099, 24'd9121410, 24'd9030702, 24'd8812923, 24'd8511174, 24'd8185169, 24'd7899424, 24'd7710487, 24'd7655750, 24'd7746043, 24'd7963499, 24'd8265083, 24'd8591112, 24'd8877066, 24'd9066355, 24'd9121519, 24'd9031641, 24'd8814508, 24'd8513090, 24'd8187037, 24'd7900875, 24'd7711234, 24'd7655644, 24'd7745106, 24'd7961916, 24'd8263167, 24'd8589243, 24'd8875614, 24'd9065606, 
24'd9121622, 24'd9032576, 24'd8816089, 24'd8515005, 24'd8188907, 24'd7902329, 24'd7711985, 24'd7655543, 24'd7744173, 24'd7960336, 24'd8261253, 24'd8587373, 24'd8874158, 24'd9064853, 24'd9121721, 24'd9033506, 24'd8817668, 24'd8516919, 24'd8190778, 24'd7903786, 24'd7712740, 24'd7655447, 24'd7743245, 24'd7958759, 24'd8259339, 24'd8585501, 24'd8872699, 24'd9064095, 24'd9121814, 24'd9034432, 
24'd8819243, 24'd8518832, 24'd8192650, 24'd7905247, 24'd7713501, 24'd7655357, 24'd7742322, 24'd7957185, 24'd8257427, 24'd8583628, 24'd8871236, 24'd9063332, 24'd9121902, 24'd9035354, 24'd8820816, 24'd8520744, 24'd8194524, 24'd7906712, 24'd7714266, 24'd7655271, 24'd7741402, 24'd7955614, 24'd8255515, 24'd8581754, 24'd8869770, 24'd9062565, 24'd9121985, 24'd9036270, 24'd8822385, 24'd8522656, 
24'd8196399, 24'd7908179, 24'd7715036, 24'd7655191, 24'd7740488, 24'd7954046, 24'd8253604, 24'd8579878, 24'd8868300, 24'd9061792, 24'd9122062, 24'd9037183, 24'd8823951, 24'd8524566, 24'd8198275, 24'd7909651, 24'd7715811, 24'd7655116, 24'd7739578, 24'd7952482, 24'd8251694, 24'd8578001, 24'd8866828, 24'd9061015, 24'd9122135, 24'd9038090, 24'd8825515, 24'd8526476, 24'd8200153, 24'd7911125, 
24'd7716590, 24'd7655046, 24'd7738672, 24'd7950920, 24'd8249785, 24'd8576123, 24'd8865352, 24'd9060234, 24'd9122202, 24'd9038994, 24'd8827075, 24'd8528384, 24'd8202032, 24'd7912603, 24'd7717374, 24'd7654981, 24'd7737771, 24'd7949361, 24'd8247877, 24'd8574243, 24'd8863872, 24'd9059447, 24'd9122264, 24'd9039892, 24'd8828632, 24'd8530292, 24'd8203912, 24'd7914084, 24'd7718163, 24'd7654921, 
24'd7736875, 24'd7947806, 24'd8245970, 24'd8572362, 24'd8862389, 24'd9058656, 24'd9122322, 24'd9040786, 24'd8830186, 24'd8532198, 24'd8205794, 24'd7915568, 24'd7718956, 24'd7654867, 24'd7735983, 24'd7946253, 24'd8244064, 24'd8570480, 24'd8860903, 24'd9057860, 24'd9122374, 24'd9041676, 24'd8831737, 24'd8534104, 24'd8207677, 24'd7917056, 24'd7719754, 24'd7654817, 24'd7735096, 24'd7944704, 
24'd8242159, 24'd8568596, 24'd8859414, 24'd9057060, 24'd9122420, 24'd9042561, 24'd8833285, 24'd8536008, 24'd8209561, 24'd7918547, 24'd7720557, 24'd7654773, 24'd7734214, 24'd7943157, 24'd8240255, 24'd8566711, 24'd8857921, 24'd9056255, 24'd9122462, 24'd9043441, 24'd8834830, 24'd8537912, 24'd8211447, 24'd7920042, 24'd7721365, 24'd7654734, 24'd7733336, 24'd7941614, 24'd8238352, 24'd8564825, 
24'd8856425, 24'd9055445, 24'd9122499, 24'd9044317, 24'd8836371, 24'd8539814, 24'd8213334, 24'd7921539, 24'd7722177, 24'd7654700, 24'd7732462, 24'd7940074, 24'd8236450, 24'd8562938, 24'd8854926, 24'd9054630, 24'd9122530, 24'd9045188, 24'd8837910, 24'd8541716, 24'd8215222, 24'd7923040, 24'd7722994, 24'd7654671, 24'd7731593, 24'd7938537, 24'd8234549, 24'd8561049, 24'd8853423, 24'd9053811, 
24'd9122556, 24'd9046054, 24'd8839445, 24'd8543616, 24'd8217111, 24'd7924544, 24'd7723815, 24'd7654648, 24'd7730729, 24'd7937003, 24'd8232649, 24'd8559159, 24'd8851917, 24'd9052987, 24'd9122577, 24'd9046916, 24'd8840977, 24'd8545515, 24'd8219001, 24'd7926052, 24'd7724642, 24'd7654629, 24'd7729869, 24'd7935473, 24'd8230751, 24'd8557268, 24'd8850408, 24'd9052158, 24'd9122593, 24'd9047774, 
24'd8842506, 24'd8547413, 24'd8220893, 24'd7927563, 24'd7725473, 24'd7654616, 24'd7729014, 24'd7933945, 24'd8228853, 24'd8555376, 24'd8848896, 24'd9051325, 24'd9122604, 24'd9048626, 24'd8844032, 24'd8549310, 24'd8222785, 24'd7929077, 24'd7726308, 24'd7654607, 24'd7728164, 24'd7932421, 24'd8226957, 24'd8553483, 24'd8847380, 24'd9050487, 24'd9122610, 24'd9049474, 24'd8845555, 24'd8551206, 
24'd8224679, 24'd7930594, 24'd7727148, 24'd7654604, 24'd7727318, 24'd7930900, 24'd8225062, 24'd8551588, 24'd8845861, 24'd9049645, 24'd9122610, 24'd9050318, 24'd8847074, 24'd8553101, 24'd8226574, 24'd7932114, 24'd7727993, 24'd7654606, 24'd7726477, 24'd7929382, 24'd8223167, 24'd8549693, 24'd8844340, 24'd9048798, 24'd9122606, 24'd9051157, 24'd8848590, 24'd8554994, 24'd8228471, 24'd7933638, 
24'd7728842, 24'd7654614, 24'd7725641, 24'd7927868, 24'd8221274, 24'd8547796, 24'd8842814, 24'd9047946, 24'd9122596, 24'd9051991, 24'd8850103, 24'd8556887, 24'd8230368, 24'd7935164, 24'd7729697, 24'd7654626, 24'd7724809, 24'd7926356, 24'd8219383, 24'd8545898, 24'd8841286, 24'd9047090, 24'd9122581, 24'd9052820, 24'd8851613, 24'd8558778, 24'd8232266, 24'd7936694, 24'd7730555, 24'd7654643, 
24'd7723982, 24'd7924848, 24'd8217492, 24'd8543999, 24'd8839754, 24'd9046229, 24'd9122561, 24'd9053645, 24'd8853120, 24'd8560668, 24'd8234166, 24'd7938227, 24'd7731419, 24'd7654666, 24'd7723159, 24'd7923343, 24'd8215603, 24'd8542099, 24'd8838220, 24'd9045363, 24'd9122536, 24'd9054465, 24'd8854623, 24'd8562557, 24'd8236066, 24'd7939764, 24'd7732286, 24'd7654694, 24'd7722341, 24'd7921842, 
24'd8213714, 24'd8540198, 24'd8836682, 24'd9044493, 24'd9122505, 24'd9055281, 24'd8856123, 24'd8564444, 24'd8237968, 24'd7941303, 24'd7733159, 24'd7654727, 24'd7721528, 24'd7920344, 24'd8211827, 24'd8538296, 24'd8835141, 24'd9043618, 24'd9122470, 24'd9056092, 24'd8857619, 24'd8566331, 24'd8239871, 24'd7942846, 24'd7734036, 24'd7654765, 24'd7720720, 24'd7918848, 24'd8209942, 24'd8536392, 
24'd8833597, 24'd9042739, 24'd9122429, 24'd9056898, 24'd8859113, 24'd8568216, 24'd8241775, 24'd7944391, 24'd7734918, 24'd7654808, 24'd7719916, 24'd7917357, 24'd8208057, 24'd8534488, 24'd8832050, 24'd9041855, 24'd9122383, 24'd9057699, 24'd8860603, 24'd8570100, 24'd8243679, 24'd7945940, 24'd7735804, 24'd7654856, 24'd7719117, 24'd7915868, 24'd8206174, 24'd8532583, 24'd8830499, 24'd9040966, 
24'd9122332, 24'd9058496, 24'd8862090, 24'd8571982, 24'd8245585, 24'd7947492, 24'd7736695, 24'd7654910, 24'd7718322, 24'd7914383, 24'd8204292, 24'd8530676, 24'd8828946, 24'd9040073, 24'd9122276, 24'd9059288, 24'd8863573, 24'd8573864, 24'd8247492, 24'd7949047, 24'd7737590, 24'd7654969, 24'd7717533, 24'd7912901, 24'd8202411, 24'd8528769, 24'd8827389, 24'd9039175, 24'd9122215, 24'd9060075, 
24'd8865053, 24'd8575744, 24'd8249400, 24'd7950605, 24'd7738490, 24'd7655032, 24'd7716748, 24'd7911423, 24'd8200532, 24'd8526861, 24'd8825830, 24'd9038273, 24'd9122149, 24'd9060858, 24'd8866530, 24'd8577622, 24'd8251309, 24'd7952166, 24'd7739395, 24'd7655101, 24'd7715967, 24'd7909948, 24'd8198654, 24'd8524952, 24'd8824267, 24'd9037366, 24'd9122077, 24'd9061636, 24'd8868004, 24'd8579500, 
24'd8253218, 24'd7953730, 24'd7740304, 24'd7655175, 24'd7715192, 24'd7908476, 24'd8196777, 24'd8523041, 24'd8822701, 24'd9036455, 24'd9122001, 24'd9062409, 24'd8869474, 24'd8581376, 24'd8255129, 24'd7955298, 24'd7741218, 24'd7655255, 24'd7714421, 24'd7907008, 24'd8194902, 24'd8521130, 24'd8821133, 24'd9035539, 24'd9121919, 24'd9063178, 24'd8870940, 24'd8583250, 24'd8257041, 24'd7956868, 
24'd7742136, 24'd7655339, 24'd7713655, 24'd7905543, 24'd8193028, 24'd8519218, 24'd8819561, 24'd9034618, 24'd9121832, 24'd9063941, 24'd8872404, 24'd8585124, 24'd8258953, 24'd7958441, 24'd7743058, 24'd7655429, 24'd7712893, 24'd7904081, 24'd8191155, 24'd8517305, 24'd8817986, 24'd9033693, 24'd9121740, 24'd9064701, 24'd8873864, 24'd8586996, 24'd8260867, 24'd7960018, 24'd7743986, 24'd7655523, 
24'd7712137, 24'd7902623, 24'd8189284, 24'd8515391, 24'd8816408, 24'd9032764, 24'd9121643, 24'd9065455, 24'd8875320, 24'd8588866, 24'd8262781, 24'd7961597, 24'd7744917, 24'd7655623, 24'd7711385, 24'd7901168, 24'd8187414, 24'd8513476, 24'd8814827, 24'd9031830, 24'd9121540, 24'd9066204, 24'd8876773, 24'd8590735, 24'd8264696, 24'd7963179, 24'd7745854, 24'd7655728, 24'd7710638, 24'd7899716, 
24'd8185546, 24'd8511561, 24'd8813243, 24'd9030891, 24'd9121433, 24'd9066949, 24'd8878223, 24'd8592603, 24'd8266612, 24'd7964765, 24'd7746795, 24'd7655838, 24'd7709895, 24'd7898268, 24'd8183679, 24'd8509644, 24'd8811657, 24'd9029948, 24'd9121320, 24'd9067689, 24'd8879669, 24'd8594469, 24'd8268529, 24'd7966353, 24'd7747740, 24'd7655953, 24'd7709158, 24'd7896824, 24'd8181813, 24'd8507727, 
24'd8810067, 24'd9029001, 24'd9121202, 24'd9068424, 24'd8881112, 24'd8596334, 24'd8270447, 24'd7967944, 24'd7748690, 24'd7656074, 24'd7708425, 24'd7895383, 24'd8179949, 24'd8505809, 24'd8808474, 24'd9028049, 24'd9121079, 24'd9069155, 24'd8882552, 24'd8598197, 24'd8272366, 24'd7969538, 24'd7749644, 24'd7656199, 24'd7707697, 24'd7893945, 24'd8178086, 24'd8503889, 24'd8806878, 24'd9027092, 
24'd9120951, 24'd9069881, 24'd8883987, 24'd8600059, 24'd8274285, 24'd7971135, 24'd7750603, 24'd7656330, 24'd7706973, 24'd7892511, 24'd8176225, 24'd8501970, 24'd8805280, 24'd9026131, 24'd9120818, 24'd9070602, 24'd8885420, 24'd8601920, 24'd8276206, 24'd7972736, 24'd7751566, 24'd7656465, 24'd7706255, 24'd7891080, 24'd8174366, 24'd8500049, 24'd8803678, 24'd9025166, 24'd9120680, 24'd9071318, 
24'd8886849, 24'd8603779, 24'd8278127, 24'd7974339, 24'd7752533, 24'd7656606, 24'd7705541, 24'd7889653, 24'd8172507, 24'd8498128, 24'd8802074, 24'd9024196, 24'd9120536, 24'd9072029, 24'd8888274, 24'd8605636, 24'd8280048, 24'd7975944, 24'd7753506, 24'd7656752, 24'd7704832, 24'd7888229, 24'd8170651, 24'd8496205, 24'd8800467, 24'd9023222, 24'd9120388, 24'd9072736, 24'd8889696, 24'd8607492, 
24'd8281971, 24'd7977553, 24'd7754482, 24'd7656903, 24'd7704128, 24'd7886809, 24'd8168795, 24'd8494282, 24'd8798856, 24'd9022243, 24'd9120234, 24'd9073438, 24'd8891115, 24'd8609346, 24'd8283894, 24'd7979165, 24'd7755463, 24'd7657060, 24'd7703428, 24'd7885392, 24'd8166942, 24'd8492359, 24'd8797243, 24'd9021260, 24'd9120075, 24'd9074135, 24'd8892530, 24'd8611199, 24'd8285818, 24'd7980779, 
24'd7756449, 24'd7657221, 24'd7702734, 24'd7883979, 24'd8165090, 24'd8490434, 24'd8795627, 24'd9020272, 24'd9119911, 24'd9074827, 24'd8893941, 24'd8613051, 24'd8287743, 24'd7982397, 24'd7757439, 24'd7657388, 24'd7702044, 24'd7882570, 24'd8163239, 24'd8488509, 24'd8794008, 24'd9019280, 24'd9119742, 24'd9075514, 24'd8895349, 24'd8614900, 24'd8289669, 24'd7984017, 24'd7758433, 24'd7657559, 
24'd7701359, 24'd7881163, 24'd8161390, 24'd8486583, 24'd8792387, 24'd9018283, 24'd9119568, 24'd9076197, 24'd8896753, 24'd8616748, 24'd8291595, 24'd7985640, 24'd7759432, 24'd7657736, 24'd7700679, 24'd7879761, 24'd8159543, 24'd8484657, 24'd8790762, 24'd9017282, 24'd9119389, 24'd9076875, 24'd8898154, 24'd8618595, 24'd8293522, 24'd7987266, 24'd7760435, 24'd7657918, 24'd7700003, 24'd7878362, 
24'd8157697, 24'd8482730, 24'd8789135, 24'd9016277, 24'd9119204, 24'd9077548, 24'd8899551, 24'd8620440, 24'd8295449, 24'd7988895, 24'd7761442, 24'd7658105, 24'd7699333, 24'd7876967, 24'd8155853, 24'd8480802, 24'd8787505, 24'd9015267, 24'd9119015, 24'd9078216, 24'd8900945, 24'd8622283, 24'd8297378, 24'd7990526, 24'd7762454, 24'd7658297, 24'd7698667, 24'd7875575, 24'd8154011, 24'd8478873, 
24'd8785872, 24'd9014253, 24'd9118820, 24'd9078879, 24'd8902335, 24'd8624125, 24'd8299306, 24'd7992160, 24'd7763471, 24'd7658494, 24'd7698006, 24'd7874187, 24'd8152170, 24'd8476944, 24'd8784236, 24'd9013234, 24'd9118620, 24'd9079537, 24'd8903721, 24'd8625965, 24'd8301236, 24'd7993798, 24'd7764492, 24'd7658697, 24'd7697350, 24'd7872802, 24'd8150331, 24'd8475014, 24'd8782598, 24'd9012211, 
24'd9118415, 24'd9080191, 24'd8905104, 24'd8627803, 24'd8303166, 24'd7995437, 24'd7765517, 24'd7658904, 24'd7696699, 24'd7871421, 24'd8148493, 24'd8473084, 24'd8780957, 24'd9011184, 24'd9118205, 24'd9080840, 24'd8906483, 24'd8629640, 24'd8305097, 24'd7997080, 24'd7766546, 24'd7659117, 24'd7696053, 24'd7870044, 24'd8146658, 24'd8471153, 24'd8779313, 24'd9010152, 24'd9117990, 24'd9081484, 
24'd8907858, 24'd8631475, 24'd8307028, 24'd7998725, 24'd7767580, 24'd7659335, 24'd7695411, 24'd7868670, 24'd8144824, 24'd8469221, 24'd8777666, 24'd9009116, 24'd9117769, 24'd9082123, 24'd8909230, 24'd8633308, 24'd8308960, 24'd8000373, 24'd7768618, 24'd7659558, 24'd7694775, 24'd7867300, 24'd8142991, 24'd8467289, 24'd8776016, 24'd9008076, 24'd9117544, 24'd9082757, 24'd8910599, 24'd8635139, 
24'd8310892, 24'd8002024, 24'd7769661, 24'd7659786, 24'd7694143, 24'd7865934, 24'd8141160, 24'd8465357, 24'd8774364, 24'd9007031, 24'd9117313, 24'd9083386, 24'd8911963, 24'd8636969, 24'd8312825, 24'd8003678, 24'd7770708, 24'd7660019, 24'd7693516, 24'd7864571, 24'd8139332, 24'd8463423, 24'd8772709, 24'd9005982, 24'd9117078, 24'd9084010, 24'd8913324, 24'd8638797, 24'd8314758, 24'd8005334, 
24'd7771759, 24'd7660257, 24'd7692894, 24'd7863212, 24'd8137504, 24'd8461490, 24'd8771052, 24'd9004929, 24'd9116837, 24'd9084630, 24'd8914681, 24'd8640624, 24'd8316692, 24'd8006993, 24'd7772814, 24'd7660500, 24'd7692277, 24'd7861856, 24'd8135679, 24'd8459556, 24'd8769392, 24'd9003871, 24'd9116591, 24'd9085245, 24'd8916035, 24'd8642448, 24'd8318627, 24'd8008655, 24'd7773874, 24'd7660749, 
24'd7691665, 24'd7860505, 24'd8133855, 24'd8457621, 24'd8767729, 24'd9002809, 24'd9116340, 24'd9085854, 24'd8917385, 24'd8644271, 24'd8320562, 24'd8010319, 24'd7774938, 24'd7661002, 24'd7691058, 24'd7859157, 24'd8132033, 24'd8455686, 24'd8766063, 24'd9001743, 24'd9116084, 24'd9086459, 24'd8918731, 24'd8646092, 24'd8322497, 24'd8011986, 24'd7776007, 24'd7661261, 24'd7690455, 24'd7857813, 
24'd8130213, 24'd8453750, 24'd8764395, 24'd9000672, 24'd9115823, 24'd9087059, 24'd8920073, 24'd8647911, 24'd8324433, 24'd8013655, 24'd7777080, 24'd7661524, 24'd7689858, 24'd7856472, 24'd8128395, 24'd8451814, 24'd8762724, 24'd8999597, 24'd9115557, 24'd9087654, 24'd8921412, 24'd8649728, 24'd8326369, 24'd8015327, 24'd7778157, 24'd7661793, 24'd7689265, 24'd7855135, 24'd8126579, 24'd8449877, 
24'd8761051, 24'd8998518, 24'd9115285, 24'd9088245, 24'd8922747, 24'd8651544, 24'd8328306, 24'd8017002, 24'd7779238, 24'd7662067, 24'd7688677, 24'd7853802, 24'd8124764, 24'd8447940, 24'd8759374, 24'd8997435, 24'd9115009, 24'd9088830, 24'd8924078, 24'd8653358, 24'd8330243, 24'd8018680, 24'd7780324, 24'd7662346, 24'd7688094, 24'd7852473, 24'd8122951, 24'd8446003, 24'd8757696, 24'd8996347, 
24'd9114727, 24'd9089410, 24'd8925405, 24'd8655169, 24'd8332181, 24'd8020360, 24'd7781414, 24'd7662630, 24'd7687516, 24'd7851147, 24'd8121140, 24'd8444065, 24'd8756014, 24'd8995255, 24'd9114441, 24'd9089986, 24'd8926729, 24'd8656979, 24'd8334119, 24'd8022042, 24'd7782508, 24'd7662919, 24'd7686943, 24'd7849825, 24'd8119331, 24'd8442127, 24'd8754331, 24'd8994159, 24'd9114149, 24'd9090556, 
24'd8928049, 24'd8658787, 24'd8336058, 24'd8023727, 24'd7783606, 24'd7663214, 24'd7686375, 24'd7848507, 24'd8117524, 24'd8440188, 24'd8752644, 24'd8993058, 24'd9113852, 24'd9091122, 24'd8929365, 24'd8660594, 24'd8337996, 24'd8025415, 24'd7784709, 24'd7663513, 24'd7685812, 24'd7847193, 24'd8115719, 24'd8438249, 24'd8750955, 24'd8991953, 24'd9113550, 24'd9091683, 24'd8930678, 24'd8662398, 
24'd8339935, 24'd8027105, 24'd7785816, 24'd7663817, 24'd7685254, 24'd7845883, 24'd8113916, 24'd8436310, 24'd8749264, 24'd8990844, 24'd9113243, 24'd9092238, 24'd8931986, 24'd8664200, 24'd8341875, 24'd8028798, 24'd7786927, 24'd7664127, 24'd7684701, 24'd7844576, 24'd8112114, 24'd8434370, 24'd8747570, 24'd8989731, 24'd9112931, 24'd9092789, 24'd8933291, 24'd8666001, 24'd8343815, 24'd8030493, 
24'd7788042, 24'd7664442, 24'd7684152, 24'd7843273, 24'd8110315, 24'd8432430, 24'd8745873, 24'd8988614, 24'd9112614, 24'd9093335, 24'd8934592, 24'd8667799, 24'd8345755, 24'd8032191, 24'd7789161, 24'd7664761, 24'd7683609, 24'd7841974, 24'd8108517, 24'd8430490, 24'd8744174, 24'd8987492, 24'd9112292, 24'd9093876, 24'd8935889, 24'd8669596, 24'd8347695, 24'd8033891, 24'd7790285, 24'd7665086, 
24'd7683070, 24'd7840679, 24'd8106722, 24'd8428549, 24'd8742473, 24'd8986366, 24'd9111965, 24'd9094412, 24'd8937182, 24'd8671390, 24'd8349636, 24'd8035594, 24'd7791413, 24'd7665416, 24'd7682537, 24'd7839388, 24'd8104928, 24'd8426609, 24'd8740768, 24'd8985236, 24'd9111632, 24'd9094943, 24'd8938471, 24'd8673183, 24'd8351577, 24'd8037299, 24'd7792545, 24'd7665751, 24'd7682008, 24'd7838100, 
24'd8103137, 24'd8424668, 24'd8739062, 24'd8984102, 24'd9111295, 24'd9095469, 24'd8939757, 24'd8674973, 24'd8353518, 24'd8039007, 24'd7793682, 24'd7666091, 24'd7681484, 24'd7836817, 24'd8101347, 24'd8422726, 24'd8737353, 24'd8982964, 24'd9110953, 24'd9095990, 24'd8941039, 24'd8676762, 24'd8355460, 24'd8040717, 24'd7794822, 24'd7666436, 24'd7680966, 24'd7835537, 24'd8099560, 24'd8420785, 
24'd8735642, 24'd8981821, 24'd9110605, 24'd9096507, 24'd8942316, 24'd8678548, 24'd8357401, 24'd8042430, 24'd7795967, 24'd7666786, 24'd7680452, 24'd7834261, 24'd8097774, 24'd8418843, 24'd8733928, 24'd8980675, 24'd9110252, 24'd9097018, 24'd8943590, 24'd8680333, 24'd8359343, 24'd8044145, 24'd7797115, 24'd7667141, 24'd7679943, 24'd7832989, 24'd8095991, 24'd8416901, 24'd8732212, 24'd8979524, 
24'd9109895, 24'd9097524, 24'd8944860, 24'd8682115, 24'd8361285, 24'd8045863, 24'd7798268, 24'd7667501, 24'd7679440, 24'd7831721, 24'd8094209, 24'd8414959, 24'd8730493, 24'd8978369, 24'd9109532, 24'd9098025, 24'd8946127, 24'd8683896, 24'd8363228, 24'd8047582, 24'd7799425, 24'd7667866, 24'd7678941, 24'd7830457, 24'd8092430, 24'd8413016, 24'd8728772, 24'd8977210, 24'd9109164, 24'd9098522, 
24'd8947389, 24'd8685674, 24'd8365170, 24'd8049305, 24'd7800587, 24'd7668237, 24'd7678447, 24'd7829197, 24'd8090653, 24'd8411074, 24'd8727048, 24'd8976046, 24'd9108791, 24'd9099013, 24'd8948647, 24'd8687450, 24'd8367113, 24'd8051029, 24'd7801752, 24'd7668612, 24'd7677958, 24'd7827940, 24'd8088878, 24'd8409131, 24'd8725323, 24'd8974879, 24'd9108413, 24'd9099500, 24'd8949901, 24'd8689224, 
24'd8369056, 24'd8052756, 24'd7802921, 24'd7668992, 24'd7677474, 24'd7826688, 24'd8087104, 24'd8407188, 24'd8723594, 24'd8973707, 24'd9108030, 24'd9099981, 24'd8951152, 24'd8690996, 24'd8370999, 24'd8054486, 24'd7804095, 24'd7669378, 24'd7676995, 24'd7825439, 24'd8085333, 24'd8405245, 24'd8721864, 24'd8972532, 24'd9107642, 24'd9100457, 24'd8952398, 24'd8692766, 24'd8372942, 24'd8056217, 
24'd7805272, 24'd7669768, 24'd7676521, 24'd7824195, 24'd8083565, 24'd8403302, 24'd8720131, 24'd8971352, 24'd9107249, 24'd9100929, 24'd8953641, 24'd8694534, 24'd8374885, 24'd8057951, 24'd7806454, 24'd7670164, 24'd7676052, 24'd7822954, 24'd8081798, 24'd8401358, 24'd8718396, 24'd8970168, 24'd9106851, 24'd9101395, 24'd8954879, 24'd8696300, 24'd8376828, 24'd8059688, 24'd7807640, 24'd7670565, 
24'd7675589, 24'd7821718, 24'd8080033, 24'd8399415, 24'd8716658, 24'd8968981, 24'd9106448, 24'd9101857, 24'd8956114, 24'd8698063, 24'd8378772, 24'd8061426, 24'd7808830, 24'd7670970, 24'd7675130, 24'd7820485, 24'd8078271, 24'd8397472, 24'd8714918, 24'd8967789, 24'd9106040, 24'd9102313, 24'd8957345, 24'd8699824, 24'd8380715, 24'd8063167, 24'd7810024, 24'd7671381, 24'd7674676, 24'd7819256, 
24'd8076511, 24'd8395528, 24'd8713176, 24'd8966593, 24'd9105627, 24'd9102764, 24'd8958571, 24'd8701584, 24'd8382658, 24'd8064911, 24'd7811222, 24'd7671797, 24'd7674227, 24'd7818032, 24'd8074753, 24'd8393585, 24'd8711432, 24'd8965393, 24'd9105209, 24'd9103211, 24'd8959794, 24'd8703341, 24'd8384602, 24'd8066656, 24'd7812424, 24'd7672217, 24'd7673783, 24'd7816811, 24'd8072997, 24'd8391641, 
24'd8709685, 24'd8964189, 24'd9104786, 24'd9103652, 24'd8961013, 24'd8705095, 24'd8386546, 24'd8068404, 24'd7813630, 24'd7672643, 24'd7673344, 24'd7815595, 24'd8071243, 24'd8389698, 24'd8707936, 24'd8962981, 24'd9104357, 24'd9104089, 24'd8962227, 24'd8706848, 24'd8388489, 24'd8070154, 24'd7814840, 24'd7673074, 24'd7672910, 24'd7814382, 24'd8069492, 24'd8387754, 24'd8706185, 24'd8961768, 
24'd9103924, 24'd9104520, 24'd8963438, 24'd8708598, 24'd8390433, 24'd8071906, 24'd7816054, 24'd7673509, 24'd7672481, 24'd7813173, 24'd8067743, 24'd8385811, 24'd8704432, 24'd8960552, 24'd9103486, 24'd9104946, 24'd8964644, 24'd8710346, 24'd8392376, 24'd8073661, 24'd7817272, 24'd7673950, 24'd7672058, 24'd7811969, 24'd8065996, 24'd8383867, 24'd8702676, 24'd8959332, 24'd9103043, 24'd9105368, 
24'd8965847, 24'd8712092, 24'd8394320, 24'd8075417, 24'd7818494, 24'd7674396, 24'd7671639, 24'd7810768, 24'd8064251, 24'd8381923, 24'd8700919, 24'd8958108, 24'd9102594, 24'd9105784, 24'd8967046, 24'd8713835, 24'd8396263, 24'd8077176, 24'd7819721, 24'd7674847, 24'd7671225, 24'd7809572, 24'd8062509, 24'd8379980, 24'd8699159, 24'd8956880, 24'd9102141, 24'd9106195, 24'd8968240, 24'd8715577, 
24'd8398207, 24'd8078937, 24'd7820951, 24'd7675303, 24'd7670816, 24'd7808379, 24'd8060769, 24'd8378037, 24'd8697396, 24'd8955648, 24'd9101683, 24'd9106601, 24'd8969430, 24'd8717316, 24'd8400150, 24'd8080700, 24'd7822185, 24'd7675763, 24'd7670412, 24'd7807191, 24'd8059031, 24'd8376093, 24'd8695632, 24'd8954412, 24'd9101219, 24'd9107002, 24'd8970617, 24'd8719052, 24'd8402093, 24'd8082466, 
24'd7823423, 24'd7676229, 24'd7670014, 24'd7806007, 24'd8057295, 24'd8374150, 24'd8693866, 24'd8953171, 24'd9100751, 24'd9107399, 24'd8971799, 24'd8720787, 24'd8404037, 24'd8084233, 24'd7824665, 24'd7676700, 24'd7669620, 24'd7804827, 24'd8055562, 24'd8372207, 24'd8692097, 24'd8951927, 24'd9100278, 24'd9107790, 24'd8972977, 24'd8722519, 24'd8405980, 24'd8086003, 24'd7825911, 24'd7677176, 
24'd7669232, 24'd7803650, 24'd8053831, 24'd8370264, 24'd8690326, 24'd8950679, 24'd9099799, 24'd9108176, 24'd8974151, 24'd8724248, 24'd8407923, 24'd8087775, 24'd7827161, 24'd7677657, 24'd7668848, 24'd7802479, 24'd8052103, 24'd8368321, 24'd8688554, 24'd8949428, 24'd9099316, 24'd9108557, 24'd8975321, 24'd8725975, 24'd8409866, 24'd8089549, 24'd7828415, 24'd7678142, 24'd7668469, 24'd7801311, 
24'd8050377, 24'd8366378, 24'd8686779, 24'd8948172, 24'd9098828, 24'd9108933, 24'd8976487, 24'd8727700, 24'd8411808, 24'd8091325, 24'd7829673, 24'd7678633, 24'd7668096, 24'd7800147, 24'd8048653, 24'd8364436, 24'd8685002, 24'd8946912, 24'd9098335, 24'd9109304, 24'd8977648, 24'd8729423, 24'd8413751, 24'd8093103, 24'd7830935, 24'd7679129, 24'd7667728, 24'd7798987, 24'd8046932, 24'd8362493, 
24'd8683223, 24'd8945648, 24'd9097836, 24'd9109670, 24'd8978806, 24'd8731143, 24'd8415693, 24'd8094883, 24'd7832200, 24'd7679629, 24'd7667364, 24'd7797832, 24'd8045213, 24'd8360551, 24'd8681441, 24'd8944381, 24'd9097333, 24'd9110031, 24'd8979959, 24'd8732861, 24'd8417635, 24'd8096665, 24'd7833470, 24'd7680135, 24'd7667006, 24'd7796680, 24'd8043496, 24'd8358609, 24'd8679658, 24'd8943109, 
24'd9096825, 24'd9110386, 24'd8981109, 24'd8734576, 24'd8419577, 24'd8098449, 24'd7834743, 24'd7680646, 24'd7666653, 24'd7795533, 24'd8041782, 24'd8356667, 24'd8677873, 24'd8941834, 24'd9096312, 24'd9110737, 24'd8982254, 24'd8736289, 24'd8421519, 24'd8100236, 24'd7836020, 24'd7681161, 24'd7666305, 24'd7794390, 24'd8040070, 24'd8354725, 24'd8676086, 24'd8940554, 24'd9095794, 24'd9111083, 
24'd8983395, 24'd8738000, 24'd8423460, 24'd8102024, 24'd7837302, 24'd7681682, 24'd7665961, 24'd7793251, 24'd8038361, 24'd8352784, 24'd8674296, 24'd8939271, 24'd9095271, 24'd9111423, 24'd8984532, 24'd8739708, 24'd8425402, 24'd8103814, 24'd7838587, 24'd7682207, 24'd7665623, 24'd7792117, 24'd8036654, 24'd8350843, 24'd8672505, 24'd8937984, 24'd9094743, 24'd9111759, 24'd8985664, 24'd8741413, 
24'd8427343, 24'd8105606, 24'd7839876, 24'd7682738, 24'd7665290, 24'd7790986, 24'd8034950, 24'd8348902, 24'd8670712, 24'd8936693, 24'd9094210, 24'd9112089, 24'd8986793, 24'd8743116, 24'd8429283, 24'd8107401, 24'd7841168, 24'd7683273, 24'd7664963, 24'd7789860, 24'd8033248, 24'd8346961, 24'd8668916, 24'd8935399, 24'd9093672, 24'd9112415, 24'd8987917, 24'd8744817, 24'd8431224, 24'd8109197, 
24'd7842465, 24'd7683814, 24'd7664640, 24'd7788738, 24'd8031549, 24'd8345021, 24'd8667119, 24'd8934100, 24'd9093129, 24'd9112735, 24'd8989037, 24'd8746515, 24'd8433164, 24'd8110995, 24'd7843766, 24'd7684359, 24'd7664322, 24'd7787620, 24'd8029852, 24'd8343081, 24'd8665320, 24'd8932798, 24'd9092582, 24'd9113050, 24'd8990153, 24'd8748211, 24'd8435104, 24'd8112795, 24'd7845070, 24'd7684909, 
24'd7664009, 24'd7786506, 24'd8028157, 24'd8341141, 24'd8663519, 24'd8931492, 24'd9092029, 24'd9113360, 24'd8991264, 24'd8749904, 24'd8437043, 24'd8114598, 24'd7846378, 24'd7685464, 24'd7663702, 24'd7785396, 24'd8026466, 24'd8339202, 24'd8661716, 24'd8930182, 24'd9091471, 24'd9113665, 24'd8992372, 24'd8751594, 24'd8438983, 24'd8116402, 24'd7847690, 24'd7686025, 24'd7663399, 24'd7784291, 
24'd8024776, 24'd8337263, 24'd8659911, 24'd8928868, 24'd9090909, 24'd9113965, 24'd8993475, 24'd8753282, 24'd8440921, 24'd8118208, 24'd7849005, 24'd7686590, 24'd7663102, 24'd7783190, 24'd8023090, 24'd8335324, 24'd8658104, 24'd8927550, 24'd9090341, 24'd9114260, 24'd8994574, 24'd8754968, 24'd8442860, 24'd8120015, 24'd7850325, 24'd7687159, 24'd7662809, 24'd7782093, 24'd8021405, 24'd8333386, 
24'd8656295, 24'd8926229, 24'd9089769, 24'd9114550, 24'd8995668, 24'd8756651, 24'd8444798, 24'd8121825, 24'd7851648, 24'd7687734, 24'd7662522, 24'd7781001, 24'd8019724, 24'd8331448, 24'd8654484, 24'd8924904, 24'd9089191, 24'd9114835, 24'd8996759, 24'd8758331, 24'd8446736, 24'd8123637, 24'd7852975, 24'd7688314, 24'd7662240, 24'd7779913, 24'd8018045, 24'd8329511, 24'd8652672, 24'd8923575, 
24'd9088609, 24'd9115114, 24'd8997845, 24'd8760009, 24'd8448673, 24'd8125450, 24'd7854306, 24'd7688899, 24'd7661963, 24'd7778829, 24'd8016368, 24'd8327574, 24'd8650857, 24'd8922242, 24'd9088022, 24'd9115389, 24'd8998927, 24'd8761684, 24'd8450610, 24'd8127265, 24'd7855640, 24'd7689488, 24'd7661691, 24'd7777749, 24'd8014695, 24'd8325637, 24'd8649041, 24'd8920906, 24'd9087430, 24'd9115658, 
24'd9000004, 24'd8763356, 24'd8452546, 24'd8129083, 24'd7856979, 24'd7690083, 24'd7661424, 24'd7776673, 24'd8013023, 24'd8323701, 24'd8647223, 24'd8919566, 24'd9086833, 24'd9115922, 24'd9001078, 24'd8765026, 24'd8454482, 24'd8130901, 24'd7858320, 24'd7690682, 24'd7661162, 24'd7775602, 24'd8011355, 24'd8321765, 24'd8645403, 24'd8918222, 24'd9086231, 24'd9116182, 24'd9002147, 24'd8766693, 
24'd8456418, 24'd8132722, 24'd7859666, 24'd7691287, 24'd7660906, 24'd7774535, 24'd8009689, 24'd8319830, 24'd8643582, 24'd8916875, 24'd9085624, 24'd9116436, 24'd9003211, 24'd8768358, 24'd8458353, 24'd8134545, 24'd7861016, 24'd7691896, 24'd7660654, 24'd7773473, 24'd8008026, 24'd8317895, 24'd8641758, 24'd8915523, 24'd9085013, 24'd9116685, 24'd9004272, 24'd8770020, 24'd8460287, 24'd8136369, 
24'd7862369, 24'd7692510, 24'd7660408, 24'd7772415, 24'd8006365, 24'd8315961, 24'd8639933, 24'd8914168, 24'd9084396, 24'd9116929, 24'd9005328, 24'd8771679, 24'd8462221, 24'd8138195, 24'd7863725, 24'd7693129, 24'd7660166, 24'd7771361, 24'd8004707, 24'd8314027, 24'd8638106, 24'd8912810, 24'd9083775, 24'd9117168, 24'd9006380, 24'd8773336, 24'd8464155, 24'd8140023, 24'd7865086, 24'd7693753, 
24'd7659930, 24'd7770311, 24'd8003052, 24'd8312094, 24'd8636277, 24'd8911448, 24'd9083149, 24'd9117401, 24'd9007427, 24'd8774989, 24'd8466088, 24'd8141853, 24'd7866450, 24'd7694381, 24'd7659699, 24'd7769266, 24'd8001400, 24'd8310161, 24'd8634447, 24'd8910082, 24'd9082517, 24'd9117630, 24'd9008470, 24'd8776641, 24'd8468020, 24'd8143684, 24'd7867818, 24'd7695015, 24'd7659473, 24'd7768225, 
24'd7999750, 24'd8308229, 24'd8632615, 24'd8908712, 24'd9081881, 24'd9117853, 24'd9009509, 24'd8778289, 24'd8469952, 24'd8145517, 24'd7869189, 24'd7695653, 24'd7659252, 24'd7767188, 24'd7998103, 24'd8306297, 24'd8630781, 24'd8907339, 24'd9081241, 24'd9118072, 24'd9010543, 24'd8779935, 24'd8471883, 24'd8147352, 24'd7870564, 24'd7696297, 24'd7659036, 24'd7766156, 24'd7996458, 24'd8304366, 
24'd8628945, 24'd8905962, 24'd9080595, 24'd9118285, 24'd9011573, 24'd8781578, 24'd8473814, 24'd8149188, 24'd7871943, 24'd7696945, 24'd7658825, 24'd7765128, 24'd7994817, 24'd8302436, 24'd8627108, 24'd8904581, 24'd9079944, 24'd9118493, 24'd9012599, 24'd8783218, 24'd8475744, 24'd8151026, 24'd7873325, 24'd7697598, 24'd7658620, 24'd7764105, 24'd7993178, 24'd8300506, 24'd8625269, 24'd8903197, 
24'd9079289, 24'd9118696, 24'd9013620, 24'd8784855, 24'd8477674, 24'd8152866, 24'd7874711, 24'd7698256, 24'd7658419, 24'd7763086, 24'd7991542, 24'd8298577, 24'd8623428, 24'd8901809, 24'd9078629, 24'd9118894, 24'd9014637, 24'd8786490, 24'd8479603, 24'd8154708, 24'd7876101, 24'd7698918, 24'd7658224, 24'd7762071, 24'd7989909, 24'd8296648, 24'd8621586, 24'd8900418, 24'd9077964, 24'd9119087, 
24'd9015650, 24'd8788122, 24'd8481531, 24'd8156551, 24'd7877494, 24'd7699586, 24'd7658034, 24'd7761061, 24'd7988278, 24'd8294720, 24'd8619742, 24'd8899023, 24'd9077294, 24'd9119274, 24'd9016658, 24'd8789751, 24'd8483458, 24'd8158395, 24'd7878891, 24'd7700258, 24'd7657849, 24'd7760055, 24'd7986651, 24'd8292793, 24'd8617897, 24'd8897625, 24'd9076619, 24'd9119457, 24'd9017661, 24'd8791377, 
24'd8485385, 24'd8160242, 24'd7880291, 24'd7700935, 24'd7657669, 24'd7759053, 24'd7985026, 24'd8290866, 24'd8616050, 24'd8896223, 24'd9075939, 24'd9119634, 24'd9018661, 24'd8793000, 24'd8487312, 24'd8162090, 24'd7881695, 24'd7701617, 24'd7657494, 24'd7758056, 24'd7983404, 24'd8288940, 24'd8614201, 24'd8894817, 24'd9075255, 24'd9119807, 24'd9019655, 24'd8794621, 24'd8489237, 24'd8163939, 
24'd7883102, 24'd7702304, 24'd7657324, 24'd7757064, 24'd7981785, 24'd8287015, 24'd8612351, 24'd8893408, 24'd9074566, 24'd9119974, 24'd9020646, 24'd8796239, 24'd8491162, 24'd8165790, 24'd7884513, 24'd7702996, 24'd7657159, 24'd7756075, 24'd7980168, 24'd8285091, 24'd8610499, 24'd8891995, 24'd9073872, 24'd9120136, 24'd9021632, 24'd8797854, 24'd8493086, 24'd8167643, 24'd7885928, 24'd7703692, 
24'd7657000, 24'd7755092, 24'd7978555, 24'd8283167, 24'd8608645, 24'd8890579, 24'd9073173, 24'd9120293, 24'd9022614, 24'd8799466, 24'd8495010, 24'd8169497, 24'd7887346, 24'd7704393, 24'd7656846, 24'd7754112, 24'd7976944, 24'd8281244, 24'd8606790, 24'd8889159, 24'd9072469, 24'd9120445, 24'd9023591, 24'd8801075, 24'd8496932, 24'd8171353, 24'd7888767, 24'd7705099, 24'd7656696, 24'd7753137, 
24'd7975337, 24'd8279322, 24'd8604934, 24'd8887736, 24'd9071761, 24'd9120591, 24'd9024563, 24'd8802681, 24'd8498854, 24'd8173210, 24'd7890192, 24'd7705810, 24'd7656552, 24'd7752167, 24'd7973732, 24'd8277400, 24'd8603076, 24'd8886309, 24'd9071048, 24'd9120733, 24'd9025532, 24'd8804284, 24'd8500775, 24'd8175069, 24'd7891621, 24'd7706526, 24'd7656413, 24'd7751201, 24'd7972130, 24'd8275479, 
24'd8601216, 24'd8884879, 24'd9070330, 24'd9120869, 24'd9026495, 24'd8805885, 24'd8502696, 24'd8176929, 24'd7893053, 24'd7707246, 24'd7656280, 24'd7750239, 24'd7970531, 24'd8273559, 24'd8599355, 24'd8883445, 24'd9069607, 24'd9121000, 24'd9027455, 24'd8807482, 24'd8504615, 24'd8178791, 24'd7894488, 24'd7707971, 24'd7656151, 24'd7749282, 24'd7968935, 24'd8271640, 24'd8597493, 24'd8882008, 
24'd9068879, 24'd9121126, 24'd9028409, 24'd8809077, 24'd8506534, 24'd8180654, 24'd7895927, 24'd7708701, 24'd7656027, 24'd7748330, 24'd7967342, 24'd8269722, 24'd8595629, 24'd8880567, 24'd9068147, 24'd9121247, 24'd9029360, 24'd8810668, 24'd8508452, 24'd8182519, 24'd7897370, 24'd7709436, 24'd7655909, 24'd7747382, 24'd7965752, 24'd8267804, 24'd8593764, 24'd8879123, 24'd9067410, 24'd9121363, 
24'd9030306, 24'd8812257, 24'd8510369, 24'd8184385, 24'd7898816, 24'd7710175, 24'd7655796, 24'd7746438, 24'd7964165, 24'd8265888, 24'd8591897, 24'd8877675, 24'd9066668, 24'd9121474, 24'd9031247, 24'd8813843, 24'd8512285, 24'd8186252, 24'd7900265, 24'd7710920, 24'd7655688, 24'd7745499, 24'd7962581, 24'd8263972, 24'd8590028, 24'd8876224, 24'd9065921, 24'd9121580, 24'd9032184, 24'd8815425, 
24'd8514201, 24'd8188121, 24'd7901718, 24'd7711669, 24'd7655585, 24'd7744565, 24'd7960999, 24'd8262057, 24'd8588159, 24'd8874770, 24'd9065170, 24'd9121680, 24'd9033116, 24'd8817005, 24'd8516115, 24'd8189992, 24'd7903174, 24'd7712422, 24'd7655487, 24'd7743634, 24'd7959421, 24'd8260143, 24'd8586288, 24'd8873312, 24'd9064414, 24'd9121775, 24'd9034044, 24'd8818582, 24'd8518029, 24'd8191863, 
24'd7904633, 24'd7713181, 24'd7655394, 24'd7742709, 24'd7957846, 24'd8258230, 24'd8584415, 24'd8871851, 24'd9063653, 24'd9121865, 24'd9034967, 24'd8820156, 24'd8519941, 24'd8193736, 24'd7906096, 24'd7713944, 24'd7655307, 24'd7741788, 24'd7956274, 24'd8256318, 24'd8582541, 24'd8870386, 24'd9062888, 24'd9121950, 24'd9035886, 24'd8821726, 24'd8521853, 24'd8195611, 24'd7907562, 24'd7714712, 
24'd7655224, 24'd7740871, 24'd7954705, 24'd8254406, 24'd8580666, 24'd8868918, 24'd9062117, 24'd9122030, 24'd9036800, 24'd8823294, 24'd8523764, 24'd8197487, 24'd7909032, 24'd7715485, 24'd7655147, 24'd7739960, 24'd7953139, 24'd8252496, 24'd8578790, 24'd8867447, 24'd9061342, 24'd9122105, 24'd9037710, 24'd8824858, 24'd8525674, 24'd8199364, 24'd7910505, 24'd7716262, 24'd7655075, 24'd7739052, 
24'd7951576, 24'd8250587, 24'd8576912, 24'd8865972, 24'd9060563, 24'd9122174, 24'd9038615, 24'd8826420, 24'd8527583, 24'd8201243, 24'd7911982, 24'd7717044, 24'd7655008, 24'd7738149, 24'd7950016, 24'd8248678, 24'd8575033, 24'd8864494, 24'd9059778, 24'd9122239, 24'd9039515, 24'd8827978, 24'd8529491, 24'd8203122, 24'd7913461, 24'd7717831, 24'd7654946, 24'd7737251, 24'd7948459, 24'd8246771, 
24'd8573152, 24'd8863013, 24'd9058989, 24'd9122298, 24'd9040411, 24'd8829534, 24'd8531398, 24'd8205004, 24'd7914944, 24'd7718622, 24'd7654889, 24'd7736357, 24'd7946905, 24'd8244864, 24'd8571270, 24'd8861528, 24'd9058195, 24'd9122352, 24'd9041303, 24'd8831086, 24'd8533304, 24'd8206886, 24'd7916431, 24'd7719419, 24'd7654838, 24'd7735468, 24'd7945354, 24'd8242959, 24'd8569387, 24'd8860040, 
24'd9057397, 24'd9122401, 24'd9042190, 24'd8832635, 24'd8535208, 24'd8208770, 24'd7917921, 24'd7720219, 24'd7654791, 24'd7734584, 24'd7943806, 24'd8241054, 24'd8567503, 24'd8858548, 24'd9056593, 24'd9122445, 24'd9043072, 24'd8834181, 24'd8537112, 24'd8210655, 24'd7919414, 24'd7721025, 24'd7654750, 24'd7733704, 24'd7942262, 24'd8239151, 24'd8565617, 24'd8857054, 24'd9055785, 24'd9122484, 
24'd9043949, 24'd8835724, 24'd8539015, 24'd8212541, 24'd7920910, 24'd7721835, 24'd7654714, 24'd7732828, 24'd7940721, 24'd8237249, 24'd8563731, 24'd8855556, 24'd9054973, 24'd9122517, 24'd9044823, 24'd8837264, 24'd8540917, 24'd8214428, 24'd7922409, 24'd7722650, 24'd7654683, 24'd7731958, 24'd7939182, 24'd8235347, 24'd8561843, 24'd8854055, 24'd9054156, 24'd9122546, 24'd9045691, 24'd8838801, 
24'd8542818, 24'd8216317, 24'd7923912, 24'd7723470, 24'd7654657, 24'd7731091, 24'd7937647, 24'd8233447, 24'd8559953, 24'd8852550, 24'd9053334, 24'd9122569, 24'd9046555, 24'd8840334, 24'd8544717, 24'd8218207, 24'd7925418, 24'd7724294, 24'd7654636, 24'd7730230, 24'd7936115, 24'd8231548, 24'd8558063, 24'd8851042, 24'd9052507, 24'd9122587, 24'd9047414, 24'd8841864, 24'd8546616, 24'd8220098, 
24'd7926928, 24'd7725123, 24'd7654621, 24'd7729373, 24'd7934587, 24'd8229650, 24'd8556171, 24'd8849531, 24'd9051676, 24'd9122600, 24'd9048269, 24'd8843392, 24'd8548513, 24'd8221990, 24'd7928440, 24'd7725957, 24'd7654610, 24'd7728521, 24'd7933061, 24'd8227753, 24'd8554278, 24'd8848017, 24'd9050840, 24'd9122608, 24'd9049119, 24'd8844915, 24'd8550410, 24'd8223884, 24'd7929956, 24'd7726795, 
24'd7654605, 24'd7727673, 24'd7931539, 24'd8225858, 24'd8552384, 24'd8846500, 24'd9049999, 24'd9122611, 24'd9049964, 24'd8846436, 24'd8552305, 24'd8225778, 24'd7931475, 24'd7727638, 24'd7654605, 24'd7726830, 24'd7930020, 24'd8223963, 24'd8550489, 24'd8844979, 24'd9049154, 24'd9122608, 24'd9050805, 24'd8847954, 24'd8554199, 24'd8227674, 24'd7932997, 24'd7728485, 24'd7654610, 24'd7725992, 
24'd7928504, 24'd8222069, 24'd8548593, 24'd8843455, 24'd9048304, 24'd9122601, 24'd9051641, 24'd8849468, 24'd8556092, 24'd8229571, 24'd7934523, 24'd7729337, 24'd7654620, 24'd7725158, 24'd7926991, 24'd8220177, 24'd8546695, 24'd8841928, 24'd9047450, 24'd9122588, 24'd9052472, 24'd8850979, 24'd8557984, 24'd8231469, 24'd7936051, 24'd7730194, 24'd7654635, 24'd7724329, 24'd7925481, 24'd8218286, 
24'd8544797, 24'd8840398, 24'd9046591, 24'd9122570, 24'd9053299, 24'd8852487, 24'd8559874, 24'd8233368, 24'd7937583, 24'd7731055, 24'd7654656, 24'd7723504, 24'd7923975, 24'd8216396, 24'd8542897, 24'd8838865, 24'd9045727, 24'd9122547, 24'd9054121, 24'd8853992, 24'd8561763, 24'd8235268, 24'd7939118, 24'd7731921, 24'd7654682, 24'd7722684, 24'd7922472, 24'd8214507, 24'd8540997, 24'd8837328, 
24'd9044859, 24'd9122519, 24'd9054939, 24'd8855493, 24'd8563652, 24'd8237169, 24'd7940656, 24'd7732792, 24'd7654712, 24'd7721869, 24'd7920973, 24'd8212620, 24'd8539095, 24'd8835789, 24'd9043986, 24'd9122485, 24'd9055752, 24'd8856991, 24'd8565538};
	
	reg [16:0] testCounter = 0;
	
	reg [23:0] audioInMono;
	always @ (*) begin
		//audioInMono = adc_right_out + adc_left_out;
		audioInMono = testWave[testCounter];
	end
	
	//Determine when the driver is in the middle of pulling a sample
	logic [7:0] driverReading = 8'd0;
	always @(posedge clk) begin
		if (chipselect && write) begin
			driverReading <= writedata;
		end	
	end
	
	wire sampleBeingTaken;
	assign sampleBeingTaken = driverReading[0];
	
	//Instantiate SFFT pipeline
 	wire [`SFFT_OUTPUT_WIDTH -1:0] SFFT_Out ;
 	wire SfftOutputValid;
 	wire outputReadError;
 	wire [`nFFT -1:0] output_address;
 	assign output_address = address[`nFFT +1:2];
 	wire [`SFFT_OUTPUT_WIDTH -1:0] Output_Why;
 
 	SFFT_Pipeline sfft(
	 	.clk(clk),
	 	.reset(reset),
	 	
	 	.SampleAmplitudeIn(audioInMono),
	 	.advanceSignal(advance),
	 	
	 	//Output BRAM IO
	 	.OutputBeingRead(sampleBeingTaken),
 		.outputReadError(outputReadError),
 		.output_address(output_address),
 		.SFFT_OutReal(SFFT_OUT),
	 	.OutputValid(SfftOutputValid),
	 	.Output_Why(Output_Why)
	 	);
	
	//Sample counter
	reg [`TIME_COUNTER_WIDTH -1:0] timeCounter = 0;
	always @(posedge SfftOutputValid) begin
		timeCounter <= timeCounter + 1;
	end
	
	/*
	//Instantiate hex decoders
	hex7seg h5( .a(Output_Why[23:20]),.y(HEX5) ), // left digit
		h4( .a(Output_Why[19:16]),.y(HEX4) ),
		h3( .a(Output_Why[15:12]),.y(HEX3) ),
		h2( .a(Output_Why[11:8]),.y(HEX2) ),
		h1( .a(Output_Why[7:4]),.y(HEX1) ),
		h0( .a(Output_Why[3:0]),.y(HEX0) );
	*/	
	
	//Instantiate hex decoders
	hex7seg h5( .a(adc_out_buffer[23:20]),.y(HEX5) ), // left digit
		h4( .a(adc_out_buffer[19:16]),.y(HEX4) ),
		h3( .a(adc_out_buffer[15:12]),.y(HEX3) ),
		h2( .a(adc_out_buffer[11:8]),.y(HEX2) ),
		h1( .a(adc_out_buffer[7:4]),.y(HEX1) ),
		h0( .a(adc_out_buffer[3:0]),.y(HEX0) );
	

	
	//Map timer counter output
	parameter readOutSize = 2048;
	reg [7:0] timer_buffer [3:0];
	integer i;
	always @(posedge clk) begin
		if (sampleBeingTaken == 0) begin
			//NOTE: Each 32bit word is written in reverse byte order, due to endian-ness of software. Avoids need for ntohl conversion
			
			//Counter -> address 0-3. Assuming 32 bit counter
			timer_buffer[3] <= timeCounter[31:24];
			timer_buffer[2] <= timeCounter[23:16];
			timer_buffer[1] <= timeCounter[15:8];
			timer_buffer[0] <= timeCounter[7:0];
		end
	end

	//Read handling
	always @(*) begin
		if (address < `NFFT*2) begin
			//Convert input address into subset of SFFT_Out
			//NOTE: Each 32bit word is written in reverse byte order, due to endian-ness of software. Avoids need for ntohl conversion
			if (address % 4 == 0) begin
				readdata = Output_Why[7:0];
				//readdata = 8'h11;
			end
			else if (address % 4 == 1) begin
				readdata = Output_Why[15:8];
				//readdata = 8'h22;
			end
			else if (address % 4 == 2) begin
				readdata = Output_Why[23:16];
				//readdata = 8'h33;
			end
			else if (address % 4 == 3) begin
				readdata = Output_Why[31:24];
				//readdata = 8'h44;
			end
		end
		else if (address[15:2] == `NFFT/2) begin
			//Send the timer counter
			readdata = timer_buffer[address[1:0]];
		end
		else begin
			//Send the valid byte
			readdata = {7'b0, ~outputReadError};
		end
	end
	
		
	//Sample inputs
	always @(posedge advance) begin
		counter <= counter + 1;
		//dac_left_in <= adc_left_out;
		//dac_right_in <= adc_right_out;
		
		dac_left_in <= testWave[testCounter];
		dac_right_in <= testWave[testCounter];
		if (testCounter == 17'd44000)
			testCounter <= 0;
		end
		else begin
			testCounter <= testCounter + 1;
		end
	end
	
	always @(posedge counter[12]) begin
		adc_out_buffer <= adc_left_out;
	end
	
endmodule


//Seven segment hex decoder
module hex7seg(input logic [3:0] a,
		output logic [6:0] y);

	always @ (a) begin
		case(a)
			0 : y = 7'b100_0000;
			1 : y = 7'b111_1001;
			2 : y = 7'b010_0100;
			3 : y = 7'b011_0000;
			4 : y = 7'b001_1001;
			5 : y = 7'b001_0010;
			6 : y = 7'b000_0010;
			7 : y = 7'b111_1000;
			8 : y = 7'b000_0000;
			9 : y = 7'b001_1000; 
			10 : y = 7'b000_1000;  //a
			11 : y = 7'b000_0011;  //b
			12 : y = 7'b100_0110;  //c
			13 : y = 7'b010_0001;  //d
			14 : y = 7'b000_0110;  //e
			15 : y = 7'b000_1110;  //f
			default: y = 7'b011_1111;
		endcase
	end
endmodule


//Debouncer for push buttons
module debouncer(input clk, input [3:0] buttonsIn, output logic [3:0] buttonsOut);
	logic [20:0] timer = 21'b0;
	
	always_ff @(posedge clk) begin
		timer <= timer - 21'b1;
	end
	
	always_ff @(negedge clk) begin
		if (timer == 0)
			buttonsOut <= buttonsIn;
	end

endmodule



